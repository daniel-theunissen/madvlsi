* SPICE3 file created from mag_ladder.ext - technology: sky130A

.subckt mag_ladder Iout D6 D5 D4 D3 D2 D1 D0 Vc Vg GND Vbn VDD
X0 a_2600_10200# Vg a_2600_8300# GND sky130_fd_pr__nfet_01v8 ad=13.5 pd=12 as=11.25 ps=11.5 w=9 l=2
X1 Iout Vg a_2600_2600# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=22.5 ps=23 w=9 l=2
X2 a_2600_8300# D3 a_1600_8000# GND sky130_fd_pr__nfet_01v8 ad=12.625 pd=15 as=1 ps=4 w=1 l=4
X3 VDD Vg a_2600_14000# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=22.5 ps=23 w=9 l=2
X4 a_400_4200# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=4
X5 a_1600_6100# Vc a_400_6100# GND sky130_fd_pr__nfet_01v8 ad=1 pd=4 as=3 ps=5 w=3 l=4
X6 a_1600_13700# Vc a_400_13700# GND sky130_fd_pr__nfet_01v8 ad=1 pd=4 as=3 ps=5 w=3 l=4
X7 a_2600_2600# Vg a_2600_4500# GND sky130_fd_pr__nfet_01v8 ad=11.25 pd=11.5 as=12.625 ps=15 w=9 l=2
X8 a_2600_14000# D0 a_1600_13700# GND sky130_fd_pr__nfet_01v8 ad=12.625 pd=15 as=1 ps=4 w=1 l=4
X9 VDD Vg a_2600_4500# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=13.5 ps=12 w=9 l=2
X10 a_400_6100# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=4
X11 a_2600_2600# D6 a_1600_2300# GND sky130_fd_pr__nfet_01v8 ad=20.75 pd=29 as=1 ps=4 w=1 l=4
X12 a_2600_4500# Vg a_2600_2600# GND sky130_fd_pr__nfet_01v8 ad=13.5 pd=12 as=11.25 ps=11.5 w=9 l=2
X13 a_2600_4500# Vg a_2600_6400# GND sky130_fd_pr__nfet_01v8 ad=11.25 pd=11.5 as=12.625 ps=15 w=9 l=2
X14 a_1600_8000# Vc a_400_8000# GND sky130_fd_pr__nfet_01v8 ad=1 pd=4 as=3 ps=5 w=3 l=4
X15 VDD Vg a_2600_6400# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=13.5 ps=12 w=9 l=2
X16 a_400_11800# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=4
X17 a_400_8000# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=4
X18 a_2600_6400# Vg a_2600_4500# GND sky130_fd_pr__nfet_01v8 ad=13.5 pd=12 as=11.25 ps=11.5 w=9 l=2
X19 a_2600_10200# Vg a_2600_12100# GND sky130_fd_pr__nfet_01v8 ad=11.25 pd=11.5 as=12.625 ps=15 w=9 l=2
X20 a_2600_4500# D5 a_1600_4200# GND sky130_fd_pr__nfet_01v8 ad=12.625 pd=15 as=1 ps=4 w=1 l=4
X21 VDD Vg a_2600_12100# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=13.5 ps=12 w=9 l=2
X22 a_1600_9900# Vc a_400_9900# GND sky130_fd_pr__nfet_01v8 ad=1 pd=4 as=3 ps=5 w=3 l=4
X23 Iout Vg a_2600_2600# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=22.5 ps=23 w=9 l=2
X24 a_2600_12100# Vg a_2600_10200# GND sky130_fd_pr__nfet_01v8 ad=13.5 pd=12 as=11.25 ps=11.5 w=9 l=2
X25 a_2600_6400# Vg a_2600_8300# GND sky130_fd_pr__nfet_01v8 ad=11.25 pd=11.5 as=12.625 ps=15 w=9 l=2
X26 VDD Vg a_2600_8300# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=13.5 ps=12 w=9 l=2
X27 a_1600_2300# Vc a_400_2300# GND sky130_fd_pr__nfet_01v8 ad=1 pd=4 as=3 ps=5 w=3 l=4
X28 a_400_9900# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=4
X29 a_400_13700# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=4
X30 a_2600_10200# D2 a_1600_9900# GND sky130_fd_pr__nfet_01v8 ad=12.625 pd=15 as=1 ps=4 w=1 l=4
X31 a_2600_8300# Vg a_2600_6400# GND sky130_fd_pr__nfet_01v8 ad=13.5 pd=12 as=11.25 ps=11.5 w=9 l=2
X32 a_2600_12100# Vg a_2600_14000# GND sky130_fd_pr__nfet_01v8 ad=11.25 pd=11.5 as=12.625 ps=15 w=9 l=2
X33 a_2600_6400# D4 a_1600_6100# GND sky130_fd_pr__nfet_01v8 ad=12.625 pd=15 as=1 ps=4 w=1 l=4
X34 a_400_2300# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=4
X35 a_2600_14000# Vg a_2600_12100# GND sky130_fd_pr__nfet_01v8 ad=13.5 pd=12 as=11.25 ps=11.5 w=9 l=2
X36 VDD Vg a_2600_14000# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=13.5 ps=12 w=9 l=2
X37 a_2600_8300# Vg a_2600_10200# GND sky130_fd_pr__nfet_01v8 ad=11.25 pd=11.5 as=12.625 ps=15 w=9 l=2
X38 VDD Vg a_2600_10200# GND sky130_fd_pr__nfet_01v8 ad=22.5 pd=23 as=13.5 ps=12 w=9 l=2
X39 a_1600_11800# Vc a_400_11800# GND sky130_fd_pr__nfet_01v8 ad=1 pd=4 as=3 ps=5 w=3 l=4
X40 a_1600_4200# Vc a_400_4200# GND sky130_fd_pr__nfet_01v8 ad=1 pd=4 as=3 ps=5 w=3 l=4
X41 a_2600_12100# D1 a_1600_11800# GND sky130_fd_pr__nfet_01v8 ad=12.625 pd=15 as=1 ps=4 w=1 l=4
.ends

