* SPICE3 file created from bias_gen.ext - technology: sky130A

.subckt bias_gen Vbn Vbp VDD GND
X0 VDD a_n4470_n620# a_n4470_n620# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X1 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X2 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X3 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X4 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X5 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X6 VDD a_n4470_n620# Vbp VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X7 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X8 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X9 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X10 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X11 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X12 a_n4470_n620# a_n10230_n3090# GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X13 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X14 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X15 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X16 Vbp Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X17 a_n10200_n3190# GND GND sky130_fd_pr__res_xhigh_po_0p35 l=17.5
X18 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X19 GND Vbp GND GND sky130_fd_pr__nfet_01v8 ad=5 pd=21 as=14.2 ps=62.8 w=10 l=10
X20 Vbn Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.2 ps=6.8 w=3 l=4
X21 VDD Vbp a_n10230_n3090# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X22 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X23 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X24 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X25 VDD Vbp Vbn VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X26 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X27 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
X28 a_n10230_n3090# a_n10230_n3090# a_n10200_n3190# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=1.5 ps=7 w=3 l=4
.ends

