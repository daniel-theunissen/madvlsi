magic
tech sky130A
timestamp 1762133376
<< polycont >>
rect -2000 1350 -1900 1400
<< locali >>
rect -50 11700 10500 11800
rect -50 11450 50 11700
rect -50 11300 150 11450
rect -1200 11240 120 11250
rect -1200 11110 -1190 11240
rect -1110 11110 120 11240
rect -1200 11100 120 11110
rect 8150 9250 9650 9400
rect -6700 9050 150 9250
rect -6700 8100 150 8300
rect -6700 7150 150 7350
rect -6700 6200 150 6400
rect -6700 5250 150 5450
rect -6700 4300 150 4500
rect -6700 3350 150 3550
rect -1100 3240 100 3250
rect -1100 3160 -1090 3240
rect -1020 3160 100 3240
rect -1100 3150 100 3160
rect 50 1650 100 3150
rect 4250 2200 4450 2350
rect 8200 2300 8500 2450
rect 4350 2100 4450 2200
rect -2250 1600 100 1650
rect -2050 1350 -2000 1400
rect -1900 1350 -1850 1400
rect -6750 540 -3250 550
rect -6750 410 -3390 540
rect -3260 410 -3250 540
rect -6750 400 -3250 410
rect -2000 50 -1900 1350
rect 4400 200 4450 600
rect 6250 540 6450 600
rect 6250 410 6260 540
rect 6440 410 6450 540
rect 6250 400 6450 410
rect 8450 200 8500 2300
rect 4400 150 8500 200
rect 8650 50 8700 9250
rect 9400 8100 9650 9250
rect 10400 8050 10500 11700
rect 10300 8000 10500 8050
rect -2000 0 8700 50
<< viali >>
rect -1190 11110 -1110 11240
rect 2450 11000 2550 11350
rect -1090 3160 -1020 3240
rect -3390 410 -3260 540
rect 6260 410 6440 540
<< metal1 >>
rect 2400 11350 2600 11400
rect -1200 11240 -1100 11250
rect -1200 11110 -1190 11240
rect -1110 11110 -1100 11240
rect -1200 3500 -1100 11110
rect 2400 11000 2450 11350
rect 2550 11000 2600 11350
rect 2400 10750 2600 11000
rect 4200 10000 4750 10900
rect 4500 9200 4750 10000
rect 4500 8400 4900 9200
rect 8150 8400 10900 9200
rect 10550 7950 10900 8400
rect 10250 7650 10900 7950
rect -1200 3240 -1000 3500
rect 8800 3300 9050 4600
rect -1200 3160 -1090 3240
rect -1020 3160 -1000 3240
rect -1200 3150 -1000 3160
rect -6700 2100 -6550 3150
rect 50 3100 150 3300
rect 0 2400 150 3100
rect 4250 2500 4950 3300
rect 8150 2500 9050 3300
rect 0 2200 50 2400
rect -6700 900 -6550 1950
rect 2700 1300 3250 2500
rect 10550 2050 10900 7650
rect 8250 1350 10900 2050
rect -4500 350 -3750 950
rect 2700 600 4450 1300
rect -3400 540 6450 550
rect -3400 410 -3390 540
rect -3260 410 6260 540
rect 6440 410 6450 540
rect -3400 400 6450 410
rect 10550 350 10900 1350
rect -4500 -200 10900 350
use bias_gen  bias_gen_0
timestamp 1762058210
transform 1 0 -1535 0 -1 1205
box -5115 -1910 1585 355
use mag_cascode_bias  mag_cascode_bias_0
timestamp 1762129613
transform -1 0 9800 0 1 4400
box -550 -250 1000 3750
use mag_current_div  mag_current_div_0
timestamp 1762129267
transform 1 0 8250 0 1 2300
box -3350 0 -50 7100
use mag_ladder  mag_ladder_0
timestamp 1762122866
transform 1 0 750 0 1 2800
box -650 -600 3550 8850
use mirror  mirror_0
timestamp 1762042913
transform 1 0 4935 0 1 1015
box -535 -465 3365 1140
<< labels >>
rlabel locali -6700 9150 -6700 9150 7 D0
port 1 w
rlabel locali -6700 8200 -6700 8200 7 D1
port 2 w
rlabel locali -6700 7250 -6700 7250 7 D2
port 3 w
rlabel locali -6700 6300 -6700 6300 7 D3
port 4 w
rlabel locali -6700 5350 -6700 5350 7 D4
port 5 w
rlabel locali -6700 4400 -6700 4400 7 D5
port 6 w
rlabel locali -6700 3450 -6700 3450 7 D6
port 7 w
rlabel metal1 -6700 2650 -6700 2650 7 VDD
port 8 w
rlabel metal1 -6700 1450 -6700 1450 7 GND
port 9 w
rlabel locali -6750 450 -6750 450 7 Iout
port 10 w
<< end >>
