magic
tech sky130A
timestamp 1762129267
<< nwell >>
rect -3300 750 -100 6950
<< nmos >>
rect -2100 350 -1800 650
rect -1600 350 -1300 650
<< pmos >>
rect -2850 6400 -2450 6700
rect -2200 6400 -1800 6700
rect -1600 6400 -1200 6700
rect -950 6400 -550 6700
rect -2200 5800 -1800 6100
rect -1600 5800 -1200 6100
rect -2850 5200 -2450 5500
rect -2200 5200 -1800 5500
rect -1600 5200 -1200 5500
rect -950 5200 -550 5500
rect -2850 4600 -2450 4900
rect -950 4600 -550 4900
rect -2850 4000 -2450 4300
rect -2200 4000 -1800 4300
rect -1600 4000 -1200 4300
rect -950 4000 -550 4300
rect -2850 3400 -2450 3700
rect -950 3400 -550 3700
rect -2850 2800 -2450 3100
rect -2200 2800 -1800 3100
rect -1600 2800 -1200 3100
rect -950 2800 -550 3100
rect -2850 2200 -2450 2500
rect -950 2200 -550 2500
rect -2850 1600 -2450 1900
rect -2200 1600 -1800 1900
rect -1600 1600 -1200 1900
rect -950 1600 -550 1900
rect -2850 1000 -2450 1300
rect -2200 1000 -1800 1300
rect -1600 1000 -1200 1300
rect -950 1000 -550 1300
<< ndiff >>
rect -2300 600 -2100 650
rect -2300 400 -2250 600
rect -2150 400 -2100 600
rect -2300 350 -2100 400
rect -1800 600 -1600 650
rect -1800 400 -1750 600
rect -1650 400 -1600 600
rect -1800 350 -1600 400
rect -1300 600 -1100 650
rect -1300 400 -1250 600
rect -1150 400 -1100 600
rect -1300 350 -1100 400
<< pdiff >>
rect -3050 6650 -2850 6700
rect -3050 6450 -3000 6650
rect -2900 6450 -2850 6650
rect -3050 6400 -2850 6450
rect -2450 6650 -2200 6700
rect -2450 6450 -2350 6650
rect -2250 6450 -2200 6650
rect -2450 6400 -2200 6450
rect -1800 6650 -1600 6700
rect -1800 6450 -1750 6650
rect -1650 6450 -1600 6650
rect -1800 6400 -1600 6450
rect -1200 6650 -950 6700
rect -1200 6450 -1150 6650
rect -1050 6450 -950 6650
rect -1200 6400 -950 6450
rect -550 6650 -350 6700
rect -550 6450 -500 6650
rect -400 6450 -350 6650
rect -550 6400 -350 6450
rect -2400 6050 -2200 6100
rect -2400 5850 -2350 6050
rect -2250 5850 -2200 6050
rect -2400 5800 -2200 5850
rect -1800 6050 -1600 6100
rect -1800 5850 -1750 6050
rect -1650 5850 -1600 6050
rect -1800 5800 -1600 5850
rect -1200 6050 -1000 6100
rect -1200 5850 -1150 6050
rect -1050 5850 -1000 6050
rect -1200 5800 -1000 5850
rect -3050 5450 -2850 5500
rect -3050 5250 -3000 5450
rect -2900 5250 -2850 5450
rect -3050 5200 -2850 5250
rect -2450 5450 -2200 5500
rect -2450 5250 -2400 5450
rect -2300 5250 -2200 5450
rect -2450 5200 -2200 5250
rect -1800 5450 -1600 5500
rect -1800 5250 -1750 5450
rect -1650 5250 -1600 5450
rect -1800 5200 -1600 5250
rect -1200 5450 -950 5500
rect -1200 5250 -1100 5450
rect -1000 5250 -950 5450
rect -1200 5200 -950 5250
rect -550 5450 -350 5500
rect -550 5250 -500 5450
rect -400 5250 -350 5450
rect -550 5200 -350 5250
rect -3050 4850 -2850 4900
rect -3050 4650 -3000 4850
rect -2900 4650 -2850 4850
rect -3050 4600 -2850 4650
rect -2450 4850 -2250 4900
rect -2450 4650 -2400 4850
rect -2300 4650 -2250 4850
rect -2450 4600 -2250 4650
rect -1150 4850 -950 4900
rect -1150 4650 -1100 4850
rect -1000 4650 -950 4850
rect -1150 4600 -950 4650
rect -550 4850 -350 4900
rect -550 4650 -500 4850
rect -400 4650 -350 4850
rect -550 4600 -350 4650
rect -3050 4250 -2850 4300
rect -3050 4050 -3000 4250
rect -2900 4050 -2850 4250
rect -3050 4000 -2850 4050
rect -2450 4250 -2200 4300
rect -2450 4050 -2400 4250
rect -2300 4050 -2200 4250
rect -2450 4000 -2200 4050
rect -1800 4250 -1600 4300
rect -1800 4050 -1750 4250
rect -1650 4050 -1600 4250
rect -1800 4000 -1600 4050
rect -1200 4250 -950 4300
rect -1200 4050 -1100 4250
rect -1000 4050 -950 4250
rect -1200 4000 -950 4050
rect -550 4250 -350 4300
rect -550 4050 -500 4250
rect -400 4050 -350 4250
rect -550 4000 -350 4050
rect -3050 3650 -2850 3700
rect -3050 3450 -3000 3650
rect -2900 3450 -2850 3650
rect -3050 3400 -2850 3450
rect -2450 3650 -2250 3700
rect -2450 3450 -2400 3650
rect -2300 3450 -2250 3650
rect -2450 3400 -2250 3450
rect -1150 3650 -950 3700
rect -1150 3450 -1100 3650
rect -1000 3450 -950 3650
rect -1150 3400 -950 3450
rect -550 3650 -350 3700
rect -550 3450 -500 3650
rect -400 3450 -350 3650
rect -550 3400 -350 3450
rect -3050 3050 -2850 3100
rect -3050 2850 -3000 3050
rect -2900 2850 -2850 3050
rect -3050 2800 -2850 2850
rect -2450 3050 -2200 3100
rect -2450 2850 -2400 3050
rect -2300 2850 -2200 3050
rect -2450 2800 -2200 2850
rect -1800 3050 -1600 3100
rect -1800 2850 -1750 3050
rect -1650 2850 -1600 3050
rect -1800 2800 -1600 2850
rect -1200 3050 -950 3100
rect -1200 2850 -1100 3050
rect -1000 2850 -950 3050
rect -1200 2800 -950 2850
rect -550 3050 -350 3100
rect -550 2850 -500 3050
rect -400 2850 -350 3050
rect -550 2800 -350 2850
rect -3050 2450 -2850 2500
rect -3050 2250 -3000 2450
rect -2900 2250 -2850 2450
rect -3050 2200 -2850 2250
rect -2450 2450 -2250 2500
rect -2450 2250 -2400 2450
rect -2300 2250 -2250 2450
rect -2450 2200 -2250 2250
rect -1150 2450 -950 2500
rect -1150 2250 -1100 2450
rect -1000 2250 -950 2450
rect -1150 2200 -950 2250
rect -550 2450 -350 2500
rect -550 2250 -500 2450
rect -400 2250 -350 2450
rect -550 2200 -350 2250
rect -3050 1850 -2850 1900
rect -3050 1650 -3000 1850
rect -2900 1650 -2850 1850
rect -3050 1600 -2850 1650
rect -2450 1850 -2200 1900
rect -2450 1650 -2350 1850
rect -2250 1650 -2200 1850
rect -2450 1600 -2200 1650
rect -1800 1850 -1600 1900
rect -1800 1650 -1750 1850
rect -1650 1650 -1600 1850
rect -1800 1600 -1600 1650
rect -1200 1850 -950 1900
rect -1200 1650 -1150 1850
rect -1050 1650 -950 1850
rect -1200 1600 -950 1650
rect -550 1850 -350 1900
rect -550 1650 -500 1850
rect -400 1650 -350 1850
rect -550 1600 -350 1650
rect -3050 1250 -2850 1300
rect -3050 1050 -3000 1250
rect -2900 1050 -2850 1250
rect -3050 1000 -2850 1050
rect -2450 1250 -2200 1300
rect -2450 1050 -2350 1250
rect -2250 1050 -2200 1250
rect -2450 1000 -2200 1050
rect -1800 1250 -1600 1300
rect -1800 1050 -1750 1250
rect -1650 1050 -1600 1250
rect -1800 1000 -1600 1050
rect -1200 1250 -950 1300
rect -1200 1050 -1150 1250
rect -1050 1050 -950 1250
rect -1200 1000 -950 1050
rect -550 1250 -350 1300
rect -550 1050 -500 1250
rect -400 1050 -350 1250
rect -550 1000 -350 1050
<< ndiffc >>
rect -2250 400 -2150 600
rect -1750 400 -1650 600
rect -1250 400 -1150 600
<< pdiffc >>
rect -3000 6450 -2900 6650
rect -2350 6450 -2250 6650
rect -1750 6450 -1650 6650
rect -1150 6450 -1050 6650
rect -500 6450 -400 6650
rect -2350 5850 -2250 6050
rect -1750 5850 -1650 6050
rect -1150 5850 -1050 6050
rect -3000 5250 -2900 5450
rect -2400 5250 -2300 5450
rect -1750 5250 -1650 5450
rect -1100 5250 -1000 5450
rect -500 5250 -400 5450
rect -3000 4650 -2900 4850
rect -2400 4650 -2300 4850
rect -1100 4650 -1000 4850
rect -500 4650 -400 4850
rect -3000 4050 -2900 4250
rect -2400 4050 -2300 4250
rect -1750 4050 -1650 4250
rect -1100 4050 -1000 4250
rect -500 4050 -400 4250
rect -3000 3450 -2900 3650
rect -2400 3450 -2300 3650
rect -1100 3450 -1000 3650
rect -500 3450 -400 3650
rect -3000 2850 -2900 3050
rect -2400 2850 -2300 3050
rect -1750 2850 -1650 3050
rect -1100 2850 -1000 3050
rect -500 2850 -400 3050
rect -3000 2250 -2900 2450
rect -2400 2250 -2300 2450
rect -1100 2250 -1000 2450
rect -500 2250 -400 2450
rect -3000 1650 -2900 1850
rect -2350 1650 -2250 1850
rect -1750 1650 -1650 1850
rect -1150 1650 -1050 1850
rect -500 1650 -400 1850
rect -3000 1050 -2900 1250
rect -2350 1050 -2250 1250
rect -1750 1050 -1650 1250
rect -1150 1050 -1050 1250
rect -500 1050 -400 1250
<< psubdiff >>
rect -2500 600 -2300 650
rect -2500 400 -2450 600
rect -2350 400 -2300 600
rect -2500 350 -2300 400
rect -1100 600 -900 650
rect -1100 400 -1050 600
rect -950 400 -900 600
rect -1100 350 -900 400
<< nsubdiff >>
rect -3250 5450 -3050 5500
rect -3250 5250 -3200 5450
rect -3100 5250 -3050 5450
rect -3250 5200 -3050 5250
rect -350 5450 -150 5500
rect -350 5250 -300 5450
rect -200 5250 -150 5450
rect -350 5200 -150 5250
rect -3250 4250 -3050 4300
rect -3250 4050 -3200 4250
rect -3100 4050 -3050 4250
rect -3250 4000 -3050 4050
rect -350 4250 -150 4300
rect -350 4050 -300 4250
rect -200 4050 -150 4250
rect -350 4000 -150 4050
rect -3250 3050 -3050 3100
rect -3250 2850 -3200 3050
rect -3100 2850 -3050 3050
rect -3250 2800 -3050 2850
rect -350 3050 -150 3100
rect -350 2850 -300 3050
rect -200 2850 -150 3050
rect -350 2800 -150 2850
rect -3250 1850 -3050 1900
rect -3250 1650 -3200 1850
rect -3100 1650 -3050 1850
rect -3250 1600 -3050 1650
rect -350 1850 -150 1900
rect -350 1650 -300 1850
rect -200 1650 -150 1850
rect -350 1600 -150 1650
<< psubdiffcont >>
rect -2450 400 -2350 600
rect -1050 400 -950 600
<< nsubdiffcont >>
rect -3200 5250 -3100 5450
rect -300 5250 -200 5450
rect -3200 4050 -3100 4250
rect -300 4050 -200 4250
rect -3200 2850 -3100 3050
rect -300 2850 -200 3050
rect -3200 1650 -3100 1850
rect -300 1650 -200 1850
<< poly >>
rect -2850 6850 -2450 6900
rect -2850 6750 -2800 6850
rect -2500 6750 -2450 6850
rect -2850 6700 -2450 6750
rect -2200 6850 -1800 6900
rect -2200 6750 -2150 6850
rect -1850 6750 -1800 6850
rect -2200 6700 -1800 6750
rect -1600 6850 -1200 6900
rect -1600 6750 -1550 6850
rect -1250 6750 -1200 6850
rect -1600 6700 -1200 6750
rect -950 6850 -550 6900
rect -950 6750 -900 6850
rect -600 6750 -550 6850
rect -950 6700 -550 6750
rect -2850 6350 -2450 6400
rect -2200 6100 -1800 6400
rect -1600 6100 -1200 6400
rect -950 6350 -550 6400
rect -2850 5500 -2450 5800
rect -2200 5500 -1800 5800
rect -1600 5500 -1200 5800
rect -950 5500 -550 5800
rect -2850 4900 -2450 5200
rect -2850 4300 -2450 4600
rect -2200 4300 -1800 5200
rect -1600 4300 -1200 5200
rect -950 4900 -550 5200
rect -950 4300 -550 4600
rect -2850 3700 -2450 4000
rect -2850 3100 -2450 3400
rect -2200 3100 -1800 4000
rect -1600 3100 -1200 4000
rect -950 3700 -550 4000
rect -950 3100 -550 3400
rect -2850 2500 -2450 2800
rect -2850 1900 -2450 2200
rect -2200 1900 -1800 2800
rect -1600 1900 -1200 2800
rect -950 2500 -550 2800
rect -950 1900 -550 2200
rect -2850 1300 -2450 1600
rect -2200 1300 -1800 1600
rect -1600 1300 -1200 1600
rect -950 1300 -550 1600
rect -2850 950 -2450 1000
rect -2850 850 -2800 950
rect -2500 850 -2450 950
rect -2850 800 -2450 850
rect -2200 950 -1800 1000
rect -2200 850 -2150 950
rect -1850 850 -1800 950
rect -2200 800 -1800 850
rect -1600 950 -1200 1000
rect -1600 850 -1550 950
rect -1250 850 -1200 950
rect -1600 800 -1200 850
rect -950 950 -550 1000
rect -950 850 -900 950
rect -600 850 -550 950
rect -950 800 -550 850
rect -2100 650 -1800 700
rect -1600 650 -1300 700
rect -2100 300 -1800 350
rect -2100 200 -2050 300
rect -1850 200 -1800 300
rect -2100 150 -1800 200
rect -1600 300 -1300 350
rect -1600 200 -1550 300
rect -1350 200 -1300 300
rect -1600 150 -1300 200
<< polycont >>
rect -2800 6750 -2500 6850
rect -2150 6750 -1850 6850
rect -1550 6750 -1250 6850
rect -900 6750 -600 6850
rect -2800 850 -2500 950
rect -2150 850 -1850 950
rect -1550 850 -1250 950
rect -900 850 -600 950
rect -2050 200 -1850 300
rect -1550 200 -1350 300
<< locali >>
rect -2850 6950 -50 7100
rect -2850 6850 -2450 6950
rect -950 6850 -550 6950
rect -2850 6750 -2800 6850
rect -2500 6750 -2450 6850
rect -2200 6750 -2150 6850
rect -1850 6750 -1550 6850
rect -1250 6750 -1200 6850
rect -950 6750 -900 6850
rect -600 6750 -550 6850
rect -1750 6700 -1650 6750
rect -3050 6650 -2850 6700
rect -3050 6450 -3000 6650
rect -2900 6450 -2850 6650
rect -3050 6400 -2850 6450
rect -2400 6650 -2200 6700
rect -2400 6450 -2350 6650
rect -2250 6450 -2200 6650
rect -2400 6050 -2200 6450
rect -2400 5850 -2350 6050
rect -2250 5850 -2200 6050
rect -2400 5800 -2200 5850
rect -1800 6650 -1600 6700
rect -1800 6450 -1750 6650
rect -1650 6450 -1600 6650
rect -1800 6050 -1600 6450
rect -1800 5850 -1750 6050
rect -1650 5850 -1600 6050
rect -1800 5800 -1600 5850
rect -1200 6650 -1000 6700
rect -1200 6450 -1150 6650
rect -1050 6450 -1000 6650
rect -1200 6050 -1000 6450
rect -550 6650 -350 6700
rect -550 6450 -500 6650
rect -400 6450 -350 6650
rect -550 6400 -350 6450
rect -1200 5850 -1150 6050
rect -1050 5850 -1000 6050
rect -1200 5800 -1000 5850
rect -2400 5750 -2250 5800
rect -3050 5550 -2250 5750
rect -3200 5450 -3100 5500
rect -3200 5200 -3100 5250
rect -3050 5450 -2850 5550
rect -1750 5500 -1650 5800
rect -1150 5750 -1000 5800
rect -1150 5550 -350 5750
rect -3050 5250 -3000 5450
rect -2900 5250 -2850 5450
rect -3050 4850 -2850 5250
rect -3050 4650 -3000 4850
rect -2900 4650 -2850 4850
rect -3050 4600 -2850 4650
rect -2450 5450 -2250 5500
rect -2450 5250 -2400 5450
rect -2300 5250 -2250 5450
rect -2450 4850 -2250 5250
rect -1800 5450 -1600 5500
rect -1800 5250 -1750 5450
rect -1650 5250 -1600 5450
rect -1800 5200 -1600 5250
rect -1150 5450 -950 5500
rect -1150 5250 -1100 5450
rect -1000 5250 -950 5450
rect -2450 4650 -2400 4850
rect -2300 4650 -2250 4850
rect -2450 4550 -2250 4650
rect -3050 4350 -2250 4550
rect -3200 4250 -3100 4300
rect -3200 4000 -3100 4050
rect -3050 4250 -2850 4350
rect -1750 4300 -1650 5200
rect -1150 4850 -950 5250
rect -1150 4650 -1100 4850
rect -1000 4650 -950 4850
rect -1150 4550 -950 4650
rect -550 5450 -350 5550
rect -550 5250 -500 5450
rect -400 5250 -350 5450
rect -550 4850 -350 5250
rect -300 5450 -200 5500
rect -300 5200 -200 5250
rect -550 4650 -500 4850
rect -400 4650 -350 4850
rect -550 4600 -350 4650
rect -1150 4350 -350 4550
rect -3050 4050 -3000 4250
rect -2900 4050 -2850 4250
rect -3050 3650 -2850 4050
rect -3050 3450 -3000 3650
rect -2900 3450 -2850 3650
rect -3050 3400 -2850 3450
rect -2450 4250 -2250 4300
rect -2450 4050 -2400 4250
rect -2300 4050 -2250 4250
rect -2450 3650 -2250 4050
rect -1800 4250 -1600 4300
rect -1800 4050 -1750 4250
rect -1650 4050 -1600 4250
rect -1800 4000 -1600 4050
rect -1150 4250 -950 4300
rect -1150 4050 -1100 4250
rect -1000 4050 -950 4250
rect -2450 3450 -2400 3650
rect -2300 3450 -2250 3650
rect -2450 3350 -2250 3450
rect -3050 3150 -2250 3350
rect -3200 3050 -3100 3100
rect -3200 2800 -3100 2850
rect -3050 3050 -2850 3150
rect -1750 3100 -1650 4000
rect -1150 3650 -950 4050
rect -1150 3450 -1100 3650
rect -1000 3450 -950 3650
rect -1150 3350 -950 3450
rect -550 4250 -350 4350
rect -550 4050 -500 4250
rect -400 4050 -350 4250
rect -550 3650 -350 4050
rect -300 4250 -200 4300
rect -300 4000 -200 4050
rect -550 3450 -500 3650
rect -400 3450 -350 3650
rect -550 3400 -350 3450
rect -1150 3150 -350 3350
rect -3050 2850 -3000 3050
rect -2900 2850 -2850 3050
rect -3050 2450 -2850 2850
rect -3050 2250 -3000 2450
rect -2900 2250 -2850 2450
rect -3050 2200 -2850 2250
rect -2450 3050 -2250 3100
rect -2450 2850 -2400 3050
rect -2300 2850 -2250 3050
rect -2450 2450 -2250 2850
rect -1800 3050 -1600 3100
rect -1800 2850 -1750 3050
rect -1650 2850 -1600 3050
rect -1800 2800 -1600 2850
rect -1150 3050 -950 3100
rect -1150 2850 -1100 3050
rect -1000 2850 -950 3050
rect -2450 2250 -2400 2450
rect -2300 2250 -2250 2450
rect -2450 2150 -2250 2250
rect -3050 1950 -2250 2150
rect -1150 2450 -950 2850
rect -1150 2250 -1100 2450
rect -1000 2250 -950 2450
rect -1150 2150 -950 2250
rect -550 3050 -350 3150
rect -550 2850 -500 3050
rect -400 2850 -350 3050
rect -550 2450 -350 2850
rect -300 3050 -200 3100
rect -300 2800 -200 2850
rect -550 2250 -500 2450
rect -400 2250 -350 2450
rect -550 2200 -350 2250
rect -1150 1950 -350 2150
rect -3200 1850 -3100 1900
rect -3200 1600 -3100 1650
rect -3050 1850 -2850 1950
rect -3050 1650 -3000 1850
rect -2900 1650 -2850 1850
rect -3050 1250 -2850 1650
rect -3050 1050 -3000 1250
rect -2900 1050 -2850 1250
rect -3050 1000 -2850 1050
rect -2400 1850 -2200 1900
rect -2400 1650 -2350 1850
rect -2250 1650 -2200 1850
rect -2400 1250 -2200 1650
rect -2400 1050 -2350 1250
rect -2250 1050 -2200 1250
rect -2400 1000 -2200 1050
rect -1800 1850 -1600 1900
rect -1800 1650 -1750 1850
rect -1650 1650 -1600 1850
rect -1800 1250 -1600 1650
rect -1800 1050 -1750 1250
rect -1650 1050 -1600 1250
rect -2850 850 -2800 950
rect -2500 850 -2150 950
rect -1850 850 -1840 950
rect -2500 600 -2100 650
rect -2500 400 -2450 600
rect -2350 400 -2250 600
rect -2150 400 -2100 600
rect -2500 350 -2100 400
rect -1800 600 -1600 1050
rect -1200 1850 -1000 1900
rect -1200 1650 -1150 1850
rect -1050 1650 -1000 1850
rect -1200 1250 -1000 1650
rect -1200 1050 -1150 1250
rect -1050 1050 -1000 1250
rect -1200 1000 -1000 1050
rect -550 1850 -350 1950
rect -550 1650 -500 1850
rect -400 1650 -350 1850
rect -550 1250 -350 1650
rect -300 1850 -200 1900
rect -300 1600 -200 1650
rect -550 1050 -500 1250
rect -400 1050 -350 1250
rect -550 1000 -350 1050
rect -1560 850 -1550 950
rect -1250 850 -900 950
rect -600 850 -550 950
rect -1800 400 -1750 600
rect -1650 400 -1600 600
rect -1800 350 -1600 400
rect -1300 600 -900 650
rect -1300 400 -1250 600
rect -1150 400 -1050 600
rect -950 400 -900 600
rect -1300 350 -900 400
rect -2050 300 -1350 350
rect -1850 200 -1550 300
rect -2050 150 -1350 200
rect -1800 0 -50 150
<< viali >>
rect -3000 6450 -2900 6650
rect -500 6450 -400 6650
rect -3200 5250 -3100 5450
rect -3200 4050 -3100 4250
rect -300 5250 -200 5450
rect -3200 2850 -3100 3050
rect -300 4050 -200 4250
rect -1750 2850 -1650 3050
rect -300 2850 -200 3050
rect -3200 1650 -3100 1850
rect -2800 850 -2500 950
rect -2150 850 -1850 950
rect -2450 400 -2350 600
rect -2250 400 -2150 600
rect -300 1650 -200 1850
rect -1550 850 -1250 950
rect -900 850 -600 950
rect -1250 400 -1150 600
rect -1050 400 -950 600
<< metal1 >>
rect -3350 6650 -50 6900
rect -3350 6450 -3000 6650
rect -2900 6450 -500 6650
rect -400 6450 -50 6650
rect -3350 6100 -50 6450
rect -3250 5450 -3050 6100
rect -3250 5250 -3200 5450
rect -3100 5250 -3050 5450
rect -3250 4250 -3050 5250
rect -3250 4050 -3200 4250
rect -3100 4050 -3050 4250
rect -3250 3050 -3050 4050
rect -350 5450 -150 6100
rect -350 5250 -300 5450
rect -200 5250 -150 5450
rect -350 4250 -150 5250
rect -350 4050 -300 4250
rect -200 4050 -150 4250
rect -3250 2850 -3200 3050
rect -3100 2850 -3050 3050
rect -3250 1850 -3050 2850
rect -3250 1650 -3200 1850
rect -3100 1650 -3050 1850
rect -3250 1600 -3050 1650
rect -1800 3050 -1600 3100
rect -1800 2850 -1750 3050
rect -1650 2850 -1600 3050
rect -1800 1000 -1600 2850
rect -350 3050 -150 4050
rect -350 2850 -300 3050
rect -200 2850 -150 3050
rect -350 1850 -150 2850
rect -350 1650 -300 1850
rect -200 1650 -150 1850
rect -350 1600 -150 1650
rect -3350 950 -50 1000
rect -3350 850 -2800 950
rect -2500 850 -2150 950
rect -1850 850 -1550 950
rect -1250 850 -900 950
rect -600 850 -50 950
rect -3350 600 -50 850
rect -3350 400 -2450 600
rect -2350 400 -2250 600
rect -2150 400 -1250 600
rect -1150 400 -1050 600
rect -950 400 -50 600
rect -3350 200 -50 400
rect -2100 150 -1800 200
rect -1600 150 -1300 200
<< labels >>
rlabel metal1 -100 550 -100 550 3 GND
port 4 e
rlabel locali -100 50 -100 50 3 Vbn2
port 3 e
rlabel metal1 -100 6500 -100 6500 3 VDD
port 2 e
rlabel locali -100 7000 -100 7000 3 Vbp
port 1 e
<< end >>
