magic
tech sky130A
magscale 1 2
timestamp 1762042913
<< nwell >>
rect -950 610 6610 2210
<< nmos >>
rect -730 -60 -130 540
rect -30 -60 570 540
rect 620 -60 1220 540
rect 1270 -60 1870 540
rect 3790 -60 4390 540
rect 4440 -60 5040 540
rect 5090 -60 5690 540
rect 5790 -60 6390 540
rect -840 -770 -240 -170
rect -140 -770 460 -170
rect 720 -770 1320 -170
rect 1420 -770 2020 -170
rect 3640 -770 4240 -170
rect 4340 -770 4940 -170
rect 5200 -770 5800 -170
rect 5900 -770 6500 -170
<< pmos >>
rect -780 1480 -180 2080
rect -80 1480 520 2080
rect 620 1480 1220 2080
rect 1320 1480 1920 2080
rect 2180 1480 2780 2080
rect 2880 1480 3480 2080
rect 3740 1480 4340 2080
rect 4440 1480 5040 2080
rect 5140 1480 5740 2080
rect 5840 1480 6440 2080
rect -730 690 -130 1290
rect -30 690 570 1290
rect 670 690 1270 1290
rect 1370 690 1970 1290
rect 3690 690 4290 1290
rect 4390 690 4990 1290
rect 5090 690 5690 1290
rect 5790 690 6390 1290
<< ndiff >>
rect -830 510 -730 540
rect -830 -30 -800 510
rect -760 -30 -730 510
rect -830 -60 -730 -30
rect -130 510 -30 540
rect -130 -30 -100 510
rect -60 -30 -30 510
rect -130 -60 -30 -30
rect 570 -60 620 540
rect 1220 -60 1270 540
rect 1870 510 1970 540
rect 1870 -30 1900 510
rect 1940 -30 1970 510
rect 3690 510 3790 540
rect 1870 -60 1970 -30
rect 3690 -30 3720 510
rect 3760 -30 3790 510
rect 3690 -60 3790 -30
rect 4390 -60 4440 540
rect 5040 -60 5090 540
rect 5690 510 5790 540
rect 5690 -30 5720 510
rect 5760 -30 5790 510
rect 5690 -60 5790 -30
rect 6390 510 6490 540
rect 6390 -30 6420 510
rect 6460 -30 6490 510
rect 6390 -60 6490 -30
rect -940 -200 -840 -170
rect -940 -740 -910 -200
rect -870 -740 -840 -200
rect -940 -770 -840 -740
rect -240 -200 -140 -170
rect -240 -740 -210 -200
rect -170 -740 -140 -200
rect -240 -770 -140 -740
rect 460 -200 560 -170
rect 460 -740 490 -200
rect 530 -740 560 -200
rect 460 -770 560 -740
rect 620 -200 720 -170
rect 620 -740 650 -200
rect 690 -740 720 -200
rect 620 -770 720 -740
rect 1320 -200 1420 -170
rect 1320 -740 1350 -200
rect 1390 -740 1420 -200
rect 1320 -770 1420 -740
rect 2020 -200 2120 -170
rect 2020 -740 2050 -200
rect 2090 -740 2120 -200
rect 2020 -770 2120 -740
rect 3540 -200 3640 -170
rect 3540 -740 3570 -200
rect 3610 -740 3640 -200
rect 3540 -770 3640 -740
rect 4240 -200 4340 -170
rect 4240 -740 4270 -200
rect 4310 -740 4340 -200
rect 4240 -770 4340 -740
rect 4940 -200 5040 -170
rect 4940 -740 4970 -200
rect 5010 -740 5040 -200
rect 4940 -770 5040 -740
rect 5100 -200 5200 -170
rect 5100 -740 5130 -200
rect 5170 -740 5200 -200
rect 5100 -770 5200 -740
rect 5800 -200 5900 -170
rect 5800 -740 5830 -200
rect 5870 -740 5900 -200
rect 5800 -770 5900 -740
rect 6500 -200 6600 -170
rect 6500 -740 6530 -200
rect 6570 -740 6600 -200
rect 6500 -770 6600 -740
<< pdiff >>
rect -880 2050 -780 2080
rect -880 1510 -850 2050
rect -810 1510 -780 2050
rect -880 1480 -780 1510
rect -180 2050 -80 2080
rect -180 1510 -150 2050
rect -110 1510 -80 2050
rect -180 1480 -80 1510
rect 520 2050 620 2080
rect 520 1510 550 2050
rect 590 1510 620 2050
rect 520 1480 620 1510
rect 1220 2050 1320 2080
rect 1220 1510 1250 2050
rect 1290 1510 1320 2050
rect 1220 1480 1320 1510
rect 1920 2050 2020 2080
rect 1920 1510 1950 2050
rect 1990 1510 2020 2050
rect 1920 1480 2020 1510
rect 2080 2050 2180 2080
rect 2080 1510 2110 2050
rect 2150 1510 2180 2050
rect 2080 1480 2180 1510
rect 2780 2050 2880 2080
rect 2780 1510 2810 2050
rect 2850 1510 2880 2050
rect 2780 1480 2880 1510
rect 3480 2050 3580 2080
rect 3480 1510 3510 2050
rect 3550 1510 3580 2050
rect 3480 1480 3580 1510
rect 3640 2050 3740 2080
rect 3640 1510 3670 2050
rect 3710 1510 3740 2050
rect 3640 1480 3740 1510
rect 4340 2050 4440 2080
rect 4340 1510 4370 2050
rect 4410 1510 4440 2050
rect 4340 1480 4440 1510
rect 5040 2050 5140 2080
rect 5040 1510 5070 2050
rect 5110 1510 5140 2050
rect 5040 1480 5140 1510
rect 5740 2050 5840 2080
rect 5740 1510 5770 2050
rect 5810 1510 5840 2050
rect 5740 1480 5840 1510
rect 6440 2050 6540 2080
rect 6440 1510 6470 2050
rect 6510 1510 6540 2050
rect 6440 1480 6540 1510
rect -830 1260 -730 1290
rect -830 720 -800 1260
rect -760 720 -730 1260
rect -830 690 -730 720
rect -130 1260 -30 1290
rect -130 720 -100 1260
rect -60 720 -30 1260
rect -130 690 -30 720
rect 570 1260 670 1290
rect 570 720 600 1260
rect 640 720 670 1260
rect 570 690 670 720
rect 1270 1260 1370 1290
rect 1270 720 1300 1260
rect 1340 720 1370 1260
rect 1270 690 1370 720
rect 1970 1260 2070 1290
rect 1970 720 2000 1260
rect 2040 720 2070 1260
rect 1970 690 2070 720
rect 3590 1260 3690 1290
rect 3590 720 3620 1260
rect 3660 720 3690 1260
rect 3590 690 3690 720
rect 4290 1260 4390 1290
rect 4290 720 4320 1260
rect 4360 720 4390 1260
rect 4290 690 4390 720
rect 4990 1260 5090 1290
rect 4990 720 5020 1260
rect 5060 720 5090 1260
rect 4990 690 5090 720
rect 5690 1260 5790 1290
rect 5690 720 5720 1260
rect 5760 720 5790 1260
rect 5690 690 5790 720
rect 6390 1260 6490 1290
rect 6390 720 6420 1260
rect 6460 720 6490 1260
rect 6390 690 6490 720
<< ndiffc >>
rect -800 -30 -760 510
rect -100 -30 -60 510
rect 1900 -30 1940 510
rect 3720 -30 3760 510
rect 5720 -30 5760 510
rect 6420 -30 6460 510
rect -910 -740 -870 -200
rect -210 -740 -170 -200
rect 490 -740 530 -200
rect 650 -740 690 -200
rect 1350 -740 1390 -200
rect 2050 -740 2090 -200
rect 3570 -740 3610 -200
rect 4270 -740 4310 -200
rect 4970 -740 5010 -200
rect 5130 -740 5170 -200
rect 5830 -740 5870 -200
rect 6530 -740 6570 -200
<< pdiffc >>
rect -850 1510 -810 2050
rect -150 1510 -110 2050
rect 550 1510 590 2050
rect 1250 1510 1290 2050
rect 1950 1510 1990 2050
rect 2110 1510 2150 2050
rect 2810 1510 2850 2050
rect 3510 1510 3550 2050
rect 3670 1510 3710 2050
rect 4370 1510 4410 2050
rect 5070 1510 5110 2050
rect 5770 1510 5810 2050
rect 6470 1510 6510 2050
rect -800 720 -760 1260
rect -100 720 -60 1260
rect 600 720 640 1260
rect 1300 720 1340 1260
rect 2000 720 2040 1260
rect 3620 720 3660 1260
rect 4320 720 4360 1260
rect 5020 720 5060 1260
rect 5720 720 5760 1260
rect 6420 720 6460 1260
<< psubdiff >>
rect -990 380 -890 410
rect -990 -30 -960 380
rect -920 -30 -890 380
rect -990 -60 -890 -30
rect 2030 380 2130 410
rect 2030 -30 2060 380
rect 2100 -30 2130 380
rect 2030 -60 2130 -30
rect 3530 380 3630 410
rect 3530 -30 3560 380
rect 3600 -30 3630 380
rect 3530 -60 3630 -30
rect 6550 380 6650 410
rect 6550 -30 6580 380
rect 6620 -30 6650 380
rect 6550 -60 6650 -30
<< nsubdiff >>
rect 2070 1260 2170 1290
rect 2070 720 2100 1260
rect 2140 720 2170 1260
rect 2070 690 2170 720
rect 3490 1260 3590 1290
rect 3490 720 3520 1260
rect 3560 720 3590 1260
rect 3490 690 3590 720
<< psubdiffcont >>
rect -960 -30 -920 380
rect 2060 -30 2100 380
rect 3560 -30 3600 380
rect 6580 -30 6620 380
<< nsubdiffcont >>
rect 2100 720 2140 1260
rect 3520 720 3560 1260
<< poly >>
rect -920 2180 -50 2200
rect -920 2130 -900 2180
rect -850 2170 -50 2180
rect -850 2130 -830 2170
rect -920 2110 -830 2130
rect -80 2110 -50 2170
rect 5710 2180 6580 2200
rect 5710 2170 6510 2180
rect 490 2110 650 2140
rect 5010 2110 5170 2140
rect 5710 2110 5740 2170
rect 6490 2130 6510 2170
rect 6560 2130 6580 2180
rect 6490 2110 6580 2130
rect -780 2080 -180 2110
rect -80 2080 520 2110
rect 620 2080 1220 2110
rect 1320 2080 1920 2110
rect 2180 2080 2780 2110
rect 2880 2080 3480 2110
rect 3740 2080 4340 2110
rect 4440 2080 5040 2110
rect 5140 2080 5740 2110
rect 5840 2080 6440 2110
rect -780 1450 -180 1480
rect -80 1450 520 1480
rect 620 1450 1220 1480
rect 1320 1450 1920 1480
rect 2180 1450 2780 1480
rect 2880 1450 3480 1480
rect 3740 1450 4340 1480
rect 4440 1450 5040 1480
rect 5140 1450 5740 1480
rect 5840 1450 6440 1480
rect -730 1400 -180 1450
rect 1320 1400 1350 1450
rect -730 1370 1350 1400
rect 2180 1400 2280 1450
rect -730 1320 -180 1370
rect 2180 1340 2200 1400
rect 2260 1340 2280 1400
rect 2180 1320 2280 1340
rect 3380 1400 3480 1450
rect 3380 1340 3400 1400
rect 3460 1340 3480 1400
rect 4310 1400 4340 1450
rect 5840 1400 6390 1450
rect 4310 1370 6390 1400
rect 3380 1320 3480 1340
rect 5840 1320 6390 1370
rect -730 1290 -130 1320
rect -30 1290 570 1320
rect 670 1290 1270 1320
rect 1370 1290 1970 1320
rect 3690 1290 4290 1320
rect 4390 1290 4990 1320
rect 5090 1290 5690 1320
rect 5790 1290 6390 1320
rect -730 660 -130 690
rect -30 670 570 690
rect 670 670 1270 690
rect 1370 670 1970 690
rect -30 660 1970 670
rect 3690 670 4290 690
rect 4390 670 4990 690
rect 5090 670 5690 690
rect 3690 660 5690 670
rect 5790 660 6390 690
rect -890 630 -700 660
rect 540 640 700 660
rect 1240 640 1400 660
rect 1940 630 2030 660
rect -890 530 -860 630
rect -730 540 -130 570
rect -30 540 570 570
rect 620 540 1220 570
rect 1270 540 1870 570
rect -950 510 -860 530
rect -950 460 -930 510
rect -880 460 -860 510
rect -950 440 -860 460
rect 2000 530 2030 630
rect 3630 630 3720 660
rect 4260 640 4420 660
rect 4960 640 5120 660
rect 6360 630 6550 660
rect 3630 530 3660 630
rect 3790 540 4390 570
rect 4440 540 5040 570
rect 5090 540 5690 570
rect 5790 540 6390 570
rect 2000 510 2090 530
rect 2000 460 2020 510
rect 2070 460 2090 510
rect 2000 440 2090 460
rect 3570 510 3660 530
rect 3570 460 3590 510
rect 3640 460 3660 510
rect 3570 440 3660 460
rect 6520 530 6550 630
rect 6520 510 6610 530
rect 6520 460 6540 510
rect 6590 460 6610 510
rect 6520 440 6610 460
rect -730 -80 -130 -60
rect -30 -80 570 -60
rect 620 -80 1220 -60
rect 1270 -80 1870 -60
rect -730 -140 1870 -80
rect 3790 -80 4390 -60
rect 4440 -80 5040 -60
rect 5090 -80 5690 -60
rect 5790 -80 6390 -60
rect 1980 -140 3670 -110
rect 3790 -140 6390 -80
rect -840 -150 2020 -140
rect -840 -170 -240 -150
rect -140 -170 460 -150
rect 720 -170 1320 -150
rect 1420 -170 2020 -150
rect 3640 -150 6500 -140
rect 3640 -170 4240 -150
rect 4340 -170 4940 -150
rect 5200 -170 5800 -150
rect 5900 -170 6500 -150
rect -840 -800 -240 -770
rect -140 -800 460 -770
rect 720 -800 1320 -770
rect 1420 -800 2020 -770
rect 3640 -800 4240 -770
rect 4340 -800 4940 -770
rect 5200 -800 5800 -770
rect 5900 -800 6500 -770
rect -1060 -820 -810 -800
rect -1060 -870 -1040 -820
rect -990 -830 -810 -820
rect -990 -870 -970 -830
rect -1060 -890 -970 -870
<< polycont >>
rect -900 2130 -850 2180
rect 6510 2130 6560 2180
rect 2200 1340 2260 1400
rect 3400 1340 3460 1400
rect -930 460 -880 510
rect 2020 460 2070 510
rect 3590 460 3640 510
rect 6540 460 6590 510
rect -1040 -870 -990 -820
<< locali >>
rect -1060 2250 1270 2280
rect -1060 2240 4440 2250
rect 1230 2210 4440 2240
rect -920 2180 -830 2200
rect -920 2130 -900 2180
rect -850 2130 -830 2180
rect -920 2110 -830 2130
rect -870 2050 -790 2110
rect -870 1510 -850 2050
rect -810 1510 -790 2050
rect -870 1490 -790 1510
rect -170 2050 -90 2070
rect -170 1510 -150 2050
rect -110 1510 -90 2050
rect -900 1450 -820 1490
rect -170 1450 -90 1510
rect 530 2050 610 2070
rect 530 1510 550 2050
rect 590 1510 610 2050
rect 530 1490 610 1510
rect 1230 2050 1310 2210
rect 1230 1510 1250 2050
rect 1290 1510 1310 2050
rect 1230 1490 1310 1510
rect 1850 2110 2170 2160
rect 1850 1450 1890 2110
rect 1930 2050 2010 2070
rect 1930 1510 1950 2050
rect 1990 1510 2010 2050
rect 1930 1490 2010 1510
rect 2090 2050 2170 2110
rect 3490 2110 3810 2160
rect 2090 1510 2110 2050
rect 2150 1510 2170 2050
rect 2090 1490 2170 1510
rect 2790 2050 2870 2070
rect 2790 1510 2810 2050
rect 2850 1510 2870 2050
rect -900 610 -860 1450
rect -170 1410 1890 1450
rect -120 1321 1360 1370
rect -1060 570 -860 610
rect -820 1260 -740 1280
rect -820 720 -800 1260
rect -760 720 -740 1260
rect -1060 -180 -1020 570
rect -820 530 -740 720
rect -120 1260 -40 1321
rect -120 720 -100 1260
rect -60 720 -40 1260
rect -120 700 -40 720
rect 580 1260 660 1280
rect 580 720 600 1260
rect 640 720 660 1260
rect 580 530 660 720
rect 1280 1260 1360 1321
rect 1970 1360 2010 1490
rect 2180 1400 2280 1420
rect 2180 1360 2200 1400
rect 1970 1340 2200 1360
rect 2260 1340 2280 1400
rect 1970 1320 2280 1340
rect 1280 720 1300 1260
rect 1340 720 1360 1260
rect 1280 680 1360 720
rect 1980 1260 2160 1280
rect 1980 720 2000 1260
rect 2040 720 2100 1260
rect 2140 720 2160 1260
rect 1980 700 2160 720
rect -950 510 -740 530
rect -950 460 -930 510
rect -880 490 -800 510
rect -880 460 -860 490
rect -950 440 -860 460
rect -980 380 -900 400
rect -980 -30 -960 380
rect -920 -30 -900 380
rect -980 -50 -900 -30
rect -820 -30 -800 490
rect -760 -30 -740 510
rect -820 -50 -740 -30
rect -120 510 -40 530
rect -120 -30 -100 510
rect -60 -30 -40 510
rect 580 510 2090 530
rect 580 480 1900 510
rect -120 -130 -40 -30
rect 1880 -30 1900 480
rect 1940 480 2020 510
rect 1940 -30 1960 480
rect 2000 460 2020 480
rect 2070 460 2090 510
rect 2000 440 2090 460
rect 1880 -50 1960 -30
rect 2040 380 2120 400
rect 2040 -30 2060 380
rect 2100 -30 2120 380
rect 2040 -50 2120 -30
rect -230 -180 -40 -130
rect 2200 -180 2240 1320
rect -1060 -200 -850 -180
rect -1060 -230 -910 -200
rect -930 -740 -910 -230
rect -870 -740 -850 -200
rect -930 -800 -850 -740
rect -230 -200 -150 -180
rect -230 -740 -210 -200
rect -170 -740 -150 -200
rect -230 -760 -150 -740
rect 470 -200 550 -180
rect 470 -740 490 -200
rect 530 -740 550 -200
rect 470 -800 550 -740
rect -1070 -820 -970 -800
rect -1070 -870 -1040 -820
rect -990 -870 -970 -820
rect -930 -840 550 -800
rect 630 -200 710 -180
rect 630 -740 650 -200
rect 690 -740 710 -200
rect 630 -800 710 -740
rect 1330 -200 1410 -180
rect 1330 -740 1350 -200
rect 1390 -740 1410 -200
rect 1330 -760 1410 -740
rect 2030 -200 2240 -180
rect 2030 -740 2050 -200
rect 2090 -220 2240 -200
rect 2090 -740 2110 -220
rect 2030 -800 2110 -740
rect 630 -840 2110 -800
rect -1070 -890 -970 -870
rect 2790 -930 2870 1510
rect 3490 2050 3570 2110
rect 3490 1510 3510 2050
rect 3550 1510 3570 2050
rect 3490 1490 3570 1510
rect 3650 2050 3730 2070
rect 3650 1510 3670 2050
rect 3710 1510 3730 2050
rect 3650 1490 3730 1510
rect 3380 1400 3480 1420
rect 3380 1340 3400 1400
rect 3460 1360 3480 1400
rect 3650 1360 3690 1490
rect 3770 1450 3810 2110
rect 4350 2070 4440 2210
rect 6490 2180 6580 2200
rect 6490 2130 6510 2180
rect 6560 2130 6580 2180
rect 6490 2110 6580 2130
rect 4350 2050 4430 2070
rect 4350 1510 4370 2050
rect 4410 1510 4430 2050
rect 4350 1490 4430 1510
rect 5050 2050 5130 2070
rect 5050 1510 5070 2050
rect 5110 1510 5130 2050
rect 5050 1490 5130 1510
rect 5750 2050 5830 2070
rect 5750 1510 5770 2050
rect 5810 1510 5830 2050
rect 5750 1450 5830 1510
rect 6450 2050 6530 2110
rect 6450 1510 6470 2050
rect 6510 1510 6530 2050
rect 6450 1490 6530 1510
rect 6480 1450 6560 1490
rect 3770 1410 5830 1450
rect 3460 1340 3690 1360
rect 3380 1320 3690 1340
rect 4300 1321 5780 1370
rect 3420 -180 3460 1320
rect 3500 1260 3680 1280
rect 3500 720 3520 1260
rect 3560 720 3620 1260
rect 3660 720 3680 1260
rect 3500 700 3680 720
rect 4300 1260 4380 1321
rect 4300 720 4320 1260
rect 4360 720 4380 1260
rect 4300 680 4380 720
rect 5000 1260 5080 1280
rect 5000 720 5020 1260
rect 5060 720 5080 1260
rect 5000 530 5080 720
rect 5700 1260 5780 1321
rect 5700 720 5720 1260
rect 5760 720 5780 1260
rect 5700 700 5780 720
rect 6400 1260 6480 1280
rect 6400 720 6420 1260
rect 6460 720 6480 1260
rect 6400 530 6480 720
rect 6520 610 6560 1450
rect 6520 570 6720 610
rect 3570 510 5080 530
rect 3570 460 3590 510
rect 3640 480 3720 510
rect 3640 460 3660 480
rect 3570 440 3660 460
rect 3540 380 3620 400
rect 3540 -30 3560 380
rect 3600 -30 3620 380
rect 3540 -50 3620 -30
rect 3700 -30 3720 480
rect 3760 480 5080 510
rect 5700 510 5780 530
rect 3760 -30 3780 480
rect 3700 -50 3780 -30
rect 5700 -30 5720 510
rect 5760 -30 5780 510
rect 5700 -130 5780 -30
rect 6400 510 6610 530
rect 6400 -30 6420 510
rect 6460 490 6540 510
rect 6460 -30 6480 490
rect 6520 460 6540 490
rect 6590 460 6610 510
rect 6520 440 6610 460
rect 6400 -50 6480 -30
rect 6560 380 6640 400
rect 6560 -30 6580 380
rect 6620 -30 6640 380
rect 6560 -50 6640 -30
rect 5700 -180 5890 -130
rect 6680 -180 6720 570
rect 3420 -200 3630 -180
rect 3420 -220 3570 -200
rect 3550 -740 3570 -220
rect 3610 -740 3630 -200
rect 3550 -800 3630 -740
rect 4250 -200 4330 -180
rect 4250 -740 4270 -200
rect 4310 -740 4330 -200
rect 4250 -760 4330 -740
rect 4950 -200 5030 -180
rect 4950 -740 4970 -200
rect 5010 -740 5030 -200
rect 4950 -800 5030 -740
rect 3550 -840 5030 -800
rect 5110 -200 5190 -180
rect 5110 -740 5130 -200
rect 5170 -740 5190 -200
rect 5110 -800 5190 -740
rect 5810 -200 5890 -180
rect 5810 -740 5830 -200
rect 5870 -740 5890 -200
rect 5810 -760 5890 -740
rect 6510 -200 6720 -180
rect 6510 -740 6530 -200
rect 6570 -230 6720 -200
rect 6570 -740 6590 -230
rect 6510 -800 6590 -740
rect 5110 -840 6590 -800
<< viali >>
rect 550 1510 590 2050
rect 2100 720 2140 1260
rect -960 -30 -920 380
rect -100 -30 -60 510
rect 2060 -30 2100 380
rect -210 -740 -170 -200
rect 1350 -740 1390 -200
rect 5070 1510 5110 2050
rect 3520 720 3560 1260
rect 3560 -30 3600 380
rect 5720 -30 5760 510
rect 6580 -30 6620 380
rect 4270 -740 4310 -200
rect 5830 -740 5870 -200
<< metal1 >>
rect -1060 2050 6720 2110
rect -1060 1510 550 2050
rect 590 1510 5070 2050
rect 5110 1510 6720 2050
rect -1060 1260 6720 1510
rect -1060 720 2100 1260
rect 2140 720 3520 1260
rect 3560 720 6720 1260
rect -1060 660 6720 720
rect -1070 510 6730 580
rect -1070 380 -100 510
rect -1070 -30 -960 380
rect -920 -30 -100 380
rect -60 380 5720 510
rect -60 -30 2060 380
rect 2100 -30 3560 380
rect 3600 -30 5720 380
rect 5760 380 6730 510
rect 5760 -30 6580 380
rect 6620 -30 6730 380
rect -1070 -200 6730 -30
rect -1070 -740 -210 -200
rect -170 -740 1350 -200
rect 1390 -740 4270 -200
rect 4310 -740 5830 -200
rect 5870 -740 6730 -200
rect -1070 -800 6730 -740
<< labels >>
rlabel locali -1060 2260 -1060 2260 7 Iin
port 0 w
rlabel locali 2820 -930 2820 -930 5 Iout
port 1 s
rlabel locali -1070 -840 -1070 -840 7 Vbn
port 2 w
rlabel metal1 -1060 1430 -1060 1430 7 VDD
port 3 w
rlabel metal1 -1070 -100 -1070 -100 7 GND
port 4 w
<< end >>
