magic
tech sky130A
timestamp 1762126425
<< nmos >>
rect -2850 6400 -2450 6700
rect -2200 6400 -1800 6700
rect -1200 6400 -800 6700
rect -550 6400 -150 6700
rect -2200 5800 -1800 6100
rect -1200 5800 -800 6100
rect -2850 5200 -2450 5500
rect -2200 5200 -1800 5500
rect -1200 5200 -800 5500
rect -550 5200 -150 5500
rect -2850 4600 -2450 4900
rect -550 4600 -150 4900
rect -2850 4000 -2450 4300
rect -2200 4000 -1800 4300
rect -1200 4000 -800 4300
rect -550 4000 -150 4300
rect -2850 3400 -2450 3700
rect -550 3400 -150 3700
rect -2850 2800 -2450 3100
rect -2200 2800 -1800 3100
rect -1200 2800 -800 3100
rect -550 2800 -150 3100
rect -2850 2200 -2450 2500
rect -550 2200 -150 2500
rect -2850 1600 -2450 1900
rect -2200 1600 -1800 1900
rect -1200 1600 -800 1900
rect -550 1600 -150 1900
rect -2850 1000 -2450 1300
rect -2200 1000 -1800 1300
rect -1200 1000 -800 1300
rect -550 1000 -150 1300
rect -2150 400 -1850 700
rect -1150 400 -850 700
<< ndiff >>
rect -3050 6650 -2850 6700
rect -3050 6450 -3000 6650
rect -2900 6450 -2850 6650
rect -3050 6400 -2850 6450
rect -2450 6650 -2200 6700
rect -2450 6450 -2350 6650
rect -2250 6450 -2200 6650
rect -2450 6400 -2200 6450
rect -1800 6650 -1600 6700
rect -1400 6650 -1200 6700
rect -1800 6450 -1750 6650
rect -1650 6450 -1600 6650
rect -1400 6450 -1350 6650
rect -1250 6450 -1200 6650
rect -1800 6400 -1600 6450
rect -1400 6400 -1200 6450
rect -800 6650 -550 6700
rect -800 6450 -750 6650
rect -650 6450 -550 6650
rect -800 6400 -550 6450
rect -150 6650 50 6700
rect -150 6450 -100 6650
rect 0 6450 50 6650
rect -150 6400 50 6450
rect -2400 6050 -2200 6100
rect -2400 5850 -2350 6050
rect -2250 5850 -2200 6050
rect -2400 5800 -2200 5850
rect -1800 6050 -1600 6100
rect -1800 5850 -1750 6050
rect -1650 5850 -1600 6050
rect -1800 5800 -1600 5850
rect -1400 6050 -1200 6100
rect -1400 5850 -1350 6050
rect -1250 5850 -1200 6050
rect -1400 5800 -1200 5850
rect -800 6050 -600 6100
rect -800 5850 -750 6050
rect -650 5850 -600 6050
rect -800 5800 -600 5850
rect -3050 5450 -2850 5500
rect -3050 5250 -3000 5450
rect -2900 5250 -2850 5450
rect -3050 5200 -2850 5250
rect -2450 5450 -2200 5500
rect -2450 5250 -2400 5450
rect -2300 5250 -2200 5450
rect -2450 5200 -2200 5250
rect -1800 5450 -1600 5500
rect -1400 5450 -1200 5500
rect -1800 5250 -1750 5450
rect -1650 5250 -1600 5450
rect -1400 5250 -1350 5450
rect -1250 5250 -1200 5450
rect -1800 5200 -1600 5250
rect -1400 5200 -1200 5250
rect -800 5450 -550 5500
rect -800 5250 -700 5450
rect -600 5250 -550 5450
rect -800 5200 -550 5250
rect -150 5450 50 5500
rect -150 5250 -100 5450
rect 0 5250 50 5450
rect -150 5200 50 5250
rect -3050 4850 -2850 4900
rect -3050 4650 -3000 4850
rect -2900 4650 -2850 4850
rect -3050 4600 -2850 4650
rect -2450 4850 -2250 4900
rect -2450 4650 -2400 4850
rect -2300 4650 -2250 4850
rect -2450 4600 -2250 4650
rect -750 4850 -550 4900
rect -750 4650 -700 4850
rect -600 4650 -550 4850
rect -750 4600 -550 4650
rect -150 4850 50 4900
rect -150 4650 -100 4850
rect 0 4650 50 4850
rect -150 4600 50 4650
rect -3050 4250 -2850 4300
rect -3050 4050 -3000 4250
rect -2900 4050 -2850 4250
rect -3050 4000 -2850 4050
rect -2450 4250 -2200 4300
rect -2450 4050 -2400 4250
rect -2300 4050 -2200 4250
rect -2450 4000 -2200 4050
rect -1800 4250 -1600 4300
rect -1400 4250 -1200 4300
rect -1800 4050 -1750 4250
rect -1650 4050 -1600 4250
rect -1400 4050 -1350 4250
rect -1250 4050 -1200 4250
rect -1800 4000 -1600 4050
rect -1400 4000 -1200 4050
rect -800 4250 -550 4300
rect -800 4050 -700 4250
rect -600 4050 -550 4250
rect -800 4000 -550 4050
rect -150 4250 50 4300
rect -150 4050 -100 4250
rect 0 4050 50 4250
rect -150 4000 50 4050
rect -3050 3650 -2850 3700
rect -3050 3450 -3000 3650
rect -2900 3450 -2850 3650
rect -3050 3400 -2850 3450
rect -2450 3650 -2250 3700
rect -2450 3450 -2400 3650
rect -2300 3450 -2250 3650
rect -2450 3400 -2250 3450
rect -750 3650 -550 3700
rect -750 3450 -700 3650
rect -600 3450 -550 3650
rect -750 3400 -550 3450
rect -150 3650 50 3700
rect -150 3450 -100 3650
rect 0 3450 50 3650
rect -150 3400 50 3450
rect -3050 3050 -2850 3100
rect -3050 2850 -3000 3050
rect -2900 2850 -2850 3050
rect -3050 2800 -2850 2850
rect -2450 3050 -2200 3100
rect -2450 2850 -2400 3050
rect -2300 2850 -2200 3050
rect -2450 2800 -2200 2850
rect -1800 3050 -1600 3100
rect -1400 3050 -1200 3100
rect -1800 2850 -1750 3050
rect -1650 2850 -1600 3050
rect -1400 2850 -1350 3050
rect -1250 2850 -1200 3050
rect -1800 2800 -1600 2850
rect -1400 2800 -1200 2850
rect -800 3050 -550 3100
rect -800 2850 -700 3050
rect -600 2850 -550 3050
rect -800 2800 -550 2850
rect -150 3050 50 3100
rect -150 2850 -100 3050
rect 0 2850 50 3050
rect -150 2800 50 2850
rect -3050 2450 -2850 2500
rect -3050 2250 -3000 2450
rect -2900 2250 -2850 2450
rect -3050 2200 -2850 2250
rect -2450 2450 -2250 2500
rect -2450 2250 -2400 2450
rect -2300 2250 -2250 2450
rect -2450 2200 -2250 2250
rect -750 2450 -550 2500
rect -750 2250 -700 2450
rect -600 2250 -550 2450
rect -750 2200 -550 2250
rect -150 2450 50 2500
rect -150 2250 -100 2450
rect 0 2250 50 2450
rect -150 2200 50 2250
rect -3050 1850 -2850 1900
rect -3050 1650 -3000 1850
rect -2900 1650 -2850 1850
rect -3050 1600 -2850 1650
rect -2450 1850 -2200 1900
rect -2450 1650 -2350 1850
rect -2250 1650 -2200 1850
rect -2450 1600 -2200 1650
rect -1800 1850 -1600 1900
rect -1400 1850 -1200 1900
rect -1800 1650 -1750 1850
rect -1650 1650 -1600 1850
rect -1400 1650 -1350 1850
rect -1250 1650 -1200 1850
rect -1800 1600 -1600 1650
rect -1400 1600 -1200 1650
rect -800 1850 -550 1900
rect -800 1650 -750 1850
rect -650 1650 -550 1850
rect -800 1600 -550 1650
rect -150 1850 50 1900
rect -150 1650 -100 1850
rect 0 1650 50 1850
rect -150 1600 50 1650
rect -3050 1250 -2850 1300
rect -3050 1050 -3000 1250
rect -2900 1050 -2850 1250
rect -3050 1000 -2850 1050
rect -2450 1250 -2200 1300
rect -2450 1050 -2350 1250
rect -2250 1050 -2200 1250
rect -2450 1000 -2200 1050
rect -1800 1250 -1600 1300
rect -1800 1050 -1750 1250
rect -1650 1050 -1600 1250
rect -1800 1000 -1600 1050
rect -1400 1250 -1200 1300
rect -1400 1050 -1350 1250
rect -1250 1050 -1200 1250
rect -1400 1000 -1200 1050
rect -800 1250 -550 1300
rect -800 1050 -750 1250
rect -650 1050 -550 1250
rect -800 1000 -550 1050
rect -150 1250 50 1300
rect -150 1050 -100 1250
rect 0 1050 50 1250
rect -150 1000 50 1050
rect -2350 650 -2150 700
rect -2350 450 -2300 650
rect -2200 450 -2150 650
rect -2350 400 -2150 450
rect -1850 650 -1650 700
rect -1850 450 -1800 650
rect -1700 450 -1650 650
rect -1850 400 -1650 450
rect -1350 650 -1150 700
rect -1350 450 -1300 650
rect -1200 450 -1150 650
rect -1350 400 -1150 450
rect -850 650 -650 700
rect -850 450 -800 650
rect -700 450 -650 650
rect -850 400 -650 450
<< ndiffc >>
rect -3000 6450 -2900 6650
rect -2350 6450 -2250 6650
rect -1750 6450 -1650 6650
rect -1350 6450 -1250 6650
rect -750 6450 -650 6650
rect -100 6450 0 6650
rect -2350 5850 -2250 6050
rect -1750 5850 -1650 6050
rect -1350 5850 -1250 6050
rect -750 5850 -650 6050
rect -3000 5250 -2900 5450
rect -2400 5250 -2300 5450
rect -1750 5250 -1650 5450
rect -1350 5250 -1250 5450
rect -700 5250 -600 5450
rect -100 5250 0 5450
rect -3000 4650 -2900 4850
rect -2400 4650 -2300 4850
rect -700 4650 -600 4850
rect -100 4650 0 4850
rect -3000 4050 -2900 4250
rect -2400 4050 -2300 4250
rect -1750 4050 -1650 4250
rect -1350 4050 -1250 4250
rect -700 4050 -600 4250
rect -100 4050 0 4250
rect -3000 3450 -2900 3650
rect -2400 3450 -2300 3650
rect -700 3450 -600 3650
rect -100 3450 0 3650
rect -3000 2850 -2900 3050
rect -2400 2850 -2300 3050
rect -1750 2850 -1650 3050
rect -1350 2850 -1250 3050
rect -700 2850 -600 3050
rect -100 2850 0 3050
rect -3000 2250 -2900 2450
rect -2400 2250 -2300 2450
rect -700 2250 -600 2450
rect -100 2250 0 2450
rect -3000 1650 -2900 1850
rect -2350 1650 -2250 1850
rect -1750 1650 -1650 1850
rect -1350 1650 -1250 1850
rect -750 1650 -650 1850
rect -100 1650 0 1850
rect -3000 1050 -2900 1250
rect -2350 1050 -2250 1250
rect -1750 1050 -1650 1250
rect -1350 1050 -1250 1250
rect -750 1050 -650 1250
rect -100 1050 0 1250
rect -2300 450 -2200 650
rect -1800 450 -1700 650
rect -1300 450 -1200 650
rect -800 450 -700 650
<< psubdiff >>
rect -1600 6650 -1400 6700
rect -1600 6450 -1550 6650
rect -1450 6450 -1400 6650
rect -1600 6400 -1400 6450
rect -3250 5450 -3050 5500
rect -3250 5250 -3200 5450
rect -3100 5250 -3050 5450
rect -3250 5200 -3050 5250
rect -1600 5450 -1400 5500
rect -1600 5250 -1550 5450
rect -1450 5250 -1400 5450
rect -1600 5200 -1400 5250
rect 50 5450 250 5500
rect 50 5250 100 5450
rect 200 5250 250 5450
rect 50 5200 250 5250
rect -3250 4250 -3050 4300
rect -3250 4050 -3200 4250
rect -3100 4050 -3050 4250
rect -3250 4000 -3050 4050
rect -1600 4250 -1400 4300
rect -1600 4050 -1550 4250
rect -1450 4050 -1400 4250
rect -1600 4000 -1400 4050
rect 50 4250 250 4300
rect 50 4050 100 4250
rect 200 4050 250 4250
rect 50 4000 250 4050
rect -3250 3050 -3050 3100
rect -3250 2850 -3200 3050
rect -3100 2850 -3050 3050
rect -3250 2800 -3050 2850
rect -1600 3050 -1400 3100
rect -1600 2850 -1550 3050
rect -1450 2850 -1400 3050
rect -1600 2800 -1400 2850
rect 50 3050 250 3100
rect 50 2850 100 3050
rect 200 2850 250 3050
rect 50 2800 250 2850
rect -3250 1850 -3050 1900
rect -3250 1650 -3200 1850
rect -3100 1650 -3050 1850
rect -3250 1600 -3050 1650
rect -1600 1850 -1400 1900
rect -1600 1650 -1550 1850
rect -1450 1650 -1400 1850
rect -1600 1600 -1400 1650
rect 50 1850 250 1900
rect 50 1650 100 1850
rect 200 1650 250 1850
rect 50 1600 250 1650
<< psubdiffcont >>
rect -1550 6450 -1450 6650
rect -3200 5250 -3100 5450
rect -1550 5250 -1450 5450
rect 100 5250 200 5450
rect -3200 4050 -3100 4250
rect -1550 4050 -1450 4250
rect 100 4050 200 4250
rect -3200 2850 -3100 3050
rect -1550 2850 -1450 3050
rect 100 2850 200 3050
rect -3200 1650 -3100 1850
rect -1550 1650 -1450 1850
rect 100 1650 200 1850
<< poly >>
rect -2850 6850 -2450 6900
rect -2850 6750 -2800 6850
rect -2500 6750 -2450 6850
rect -2850 6700 -2450 6750
rect -2200 6850 -1800 6900
rect -2200 6750 -2150 6850
rect -1850 6750 -1800 6850
rect -2200 6700 -1800 6750
rect -1200 6850 -800 6900
rect -1200 6750 -1150 6850
rect -850 6750 -800 6850
rect -1200 6700 -800 6750
rect -550 6850 -150 6900
rect -550 6750 -500 6850
rect -200 6750 -150 6850
rect -550 6700 -150 6750
rect -2850 6350 -2450 6400
rect -2200 6100 -1800 6400
rect -1200 6100 -800 6400
rect -550 6350 -150 6400
rect -2850 5500 -2450 5800
rect -2200 5500 -1800 5800
rect -1200 5500 -800 5800
rect -550 5500 -150 5800
rect -2850 4900 -2450 5200
rect -2850 4300 -2450 4600
rect -2200 4300 -1800 5200
rect -1200 4300 -800 5200
rect -550 4900 -150 5200
rect -550 4300 -150 4600
rect -2850 3700 -2450 4000
rect -2850 3100 -2450 3400
rect -2200 3100 -1800 4000
rect -1200 3100 -800 4000
rect -550 3700 -150 4000
rect -550 3100 -150 3400
rect -2850 2500 -2450 2800
rect -2850 1900 -2450 2200
rect -2200 1900 -1800 2800
rect -1200 1900 -800 2800
rect -550 2500 -150 2800
rect -550 1900 -150 2200
rect -2850 1300 -2450 1600
rect -2200 1300 -1800 1600
rect -1200 1300 -800 1600
rect -550 1300 -150 1600
rect -2850 950 -2450 1000
rect -2850 850 -2800 950
rect -2500 850 -2450 950
rect -2850 800 -2450 850
rect -2200 950 -1800 1000
rect -2200 850 -2150 950
rect -1850 850 -1800 950
rect -2200 800 -1800 850
rect -1200 950 -800 1000
rect -1200 850 -1150 950
rect -850 850 -800 950
rect -1200 800 -800 850
rect -550 950 -150 1000
rect -550 850 -500 950
rect -200 850 -150 950
rect -550 800 -150 850
rect -2150 700 -1850 750
rect -1150 700 -850 750
rect -2150 350 -1850 400
rect -2150 250 -2100 350
rect -1900 250 -1850 350
rect -2150 200 -1850 250
rect -1150 350 -850 400
rect -1150 250 -1100 350
rect -900 250 -850 350
rect -1150 200 -850 250
<< polycont >>
rect -2800 6750 -2500 6850
rect -2150 6750 -1850 6850
rect -1150 6750 -850 6850
rect -500 6750 -200 6850
rect -2800 850 -2500 950
rect -2150 850 -1850 950
rect -1150 850 -850 950
rect -500 850 -200 950
rect -2100 250 -1900 350
rect -1100 250 -900 350
<< locali >>
rect -2850 6950 300 7100
rect -2850 6850 -2450 6950
rect -550 6850 -150 6950
rect -2850 6750 -2800 6850
rect -2500 6750 -2450 6850
rect -2200 6750 -2150 6850
rect -1850 6750 -1150 6850
rect -850 6750 -800 6850
rect -550 6750 -500 6850
rect -200 6750 -150 6850
rect -1750 6700 -1650 6750
rect -1350 6700 -1250 6750
rect -3050 6650 -2850 6700
rect -3050 6450 -3000 6650
rect -2900 6450 -2850 6650
rect -3050 6400 -2850 6450
rect -2400 6650 -2200 6700
rect -2400 6450 -2350 6650
rect -2250 6450 -2200 6650
rect -2400 6050 -2200 6450
rect -2400 5850 -2350 6050
rect -2250 5850 -2200 6050
rect -2400 5800 -2200 5850
rect -1800 6650 -1600 6700
rect -1800 6450 -1750 6650
rect -1650 6450 -1600 6650
rect -1800 6050 -1600 6450
rect -1550 6650 -1450 6700
rect -1550 6400 -1450 6450
rect -1400 6650 -1200 6700
rect -1400 6450 -1350 6650
rect -1250 6450 -1200 6650
rect -1800 5850 -1750 6050
rect -1650 5850 -1600 6050
rect -1800 5800 -1600 5850
rect -1400 6050 -1200 6450
rect -1400 5850 -1350 6050
rect -1250 5850 -1200 6050
rect -1400 5800 -1200 5850
rect -800 6650 -600 6700
rect -800 6450 -750 6650
rect -650 6450 -600 6650
rect -800 6050 -600 6450
rect -150 6650 50 6700
rect -150 6450 -100 6650
rect 0 6450 50 6650
rect -150 6400 50 6450
rect -800 5850 -750 6050
rect -650 5850 -600 6050
rect -800 5800 -600 5850
rect -2400 5750 -2250 5800
rect -3050 5550 -2250 5750
rect -3200 5450 -3100 5500
rect -3200 5200 -3100 5250
rect -3050 5450 -2850 5550
rect -1750 5500 -1650 5800
rect -1350 5500 -1250 5800
rect -750 5750 -600 5800
rect -750 5550 50 5750
rect -3050 5250 -3000 5450
rect -2900 5250 -2850 5450
rect -3050 4850 -2850 5250
rect -3050 4650 -3000 4850
rect -2900 4650 -2850 4850
rect -3050 4600 -2850 4650
rect -2450 5450 -2250 5500
rect -2450 5250 -2400 5450
rect -2300 5250 -2250 5450
rect -2450 4850 -2250 5250
rect -1800 5450 -1600 5500
rect -1800 5250 -1750 5450
rect -1650 5250 -1600 5450
rect -1800 5200 -1600 5250
rect -1550 5450 -1450 5500
rect -1550 5200 -1450 5250
rect -1400 5450 -1200 5500
rect -1400 5250 -1350 5450
rect -1250 5250 -1200 5450
rect -1400 5200 -1200 5250
rect -750 5450 -550 5500
rect -750 5250 -700 5450
rect -600 5250 -550 5450
rect -2450 4650 -2400 4850
rect -2300 4650 -2250 4850
rect -2450 4550 -2250 4650
rect -3050 4350 -2250 4550
rect -3200 4250 -3100 4300
rect -3200 4000 -3100 4050
rect -3050 4250 -2850 4350
rect -1750 4300 -1650 5200
rect -1350 4300 -1250 5200
rect -750 4850 -550 5250
rect -750 4650 -700 4850
rect -600 4650 -550 4850
rect -750 4550 -550 4650
rect -150 5450 50 5550
rect -150 5250 -100 5450
rect 0 5250 50 5450
rect -150 4850 50 5250
rect 100 5450 200 5500
rect 100 5200 200 5250
rect -150 4650 -100 4850
rect 0 4650 50 4850
rect -150 4600 50 4650
rect -750 4350 50 4550
rect -3050 4050 -3000 4250
rect -2900 4050 -2850 4250
rect -3050 3650 -2850 4050
rect -3050 3450 -3000 3650
rect -2900 3450 -2850 3650
rect -3050 3400 -2850 3450
rect -2450 4250 -2250 4300
rect -2450 4050 -2400 4250
rect -2300 4050 -2250 4250
rect -2450 3650 -2250 4050
rect -1800 4250 -1600 4300
rect -1800 4050 -1750 4250
rect -1650 4050 -1600 4250
rect -1800 4000 -1600 4050
rect -1550 4250 -1450 4300
rect -1550 4000 -1450 4050
rect -1400 4250 -1200 4300
rect -1400 4050 -1350 4250
rect -1250 4050 -1200 4250
rect -1400 4000 -1200 4050
rect -750 4250 -550 4300
rect -750 4050 -700 4250
rect -600 4050 -550 4250
rect -2450 3450 -2400 3650
rect -2300 3450 -2250 3650
rect -2450 3350 -2250 3450
rect -3050 3150 -2250 3350
rect -3200 3050 -3100 3100
rect -3200 2800 -3100 2850
rect -3050 3050 -2850 3150
rect -1750 3100 -1650 4000
rect -1350 3100 -1250 4000
rect -750 3650 -550 4050
rect -750 3450 -700 3650
rect -600 3450 -550 3650
rect -750 3350 -550 3450
rect -150 4250 50 4350
rect -150 4050 -100 4250
rect 0 4050 50 4250
rect -150 3650 50 4050
rect 100 4250 200 4300
rect 100 4000 200 4050
rect -150 3450 -100 3650
rect 0 3450 50 3650
rect -150 3400 50 3450
rect -750 3150 50 3350
rect -3050 2850 -3000 3050
rect -2900 2850 -2850 3050
rect -3050 2450 -2850 2850
rect -3050 2250 -3000 2450
rect -2900 2250 -2850 2450
rect -3050 2200 -2850 2250
rect -2450 3050 -2250 3100
rect -2450 2850 -2400 3050
rect -2300 2850 -2250 3050
rect -2450 2450 -2250 2850
rect -1800 3050 -1600 3100
rect -1800 2850 -1750 3050
rect -1650 2850 -1600 3050
rect -1800 2800 -1600 2850
rect -1550 3050 -1450 3100
rect -1550 2800 -1450 2850
rect -1400 3050 -1200 3100
rect -1400 2850 -1350 3050
rect -1250 2850 -1200 3050
rect -1400 2800 -1200 2850
rect -750 3050 -550 3100
rect -750 2850 -700 3050
rect -600 2850 -550 3050
rect -2450 2250 -2400 2450
rect -2300 2250 -2250 2450
rect -2450 2150 -2250 2250
rect -3050 1950 -2250 2150
rect -750 2450 -550 2850
rect -750 2250 -700 2450
rect -600 2250 -550 2450
rect -750 2150 -550 2250
rect -150 3050 50 3150
rect -150 2850 -100 3050
rect 0 2850 50 3050
rect -150 2450 50 2850
rect 100 3050 200 3100
rect 100 2800 200 2850
rect -150 2250 -100 2450
rect 0 2250 50 2450
rect -150 2200 50 2250
rect -750 1950 50 2150
rect -3200 1850 -3100 1900
rect -3200 1600 -3100 1650
rect -3050 1850 -2850 1950
rect -3050 1650 -3000 1850
rect -2900 1650 -2850 1850
rect -3050 1250 -2850 1650
rect -3050 1050 -3000 1250
rect -2900 1050 -2850 1250
rect -3050 1000 -2850 1050
rect -2400 1850 -2200 1900
rect -2400 1650 -2350 1850
rect -2250 1650 -2200 1850
rect -2400 1250 -2200 1650
rect -2400 1050 -2350 1250
rect -2250 1050 -2200 1250
rect -2400 1000 -2200 1050
rect -1800 1850 -1600 1900
rect -1800 1650 -1750 1850
rect -1650 1650 -1600 1850
rect -1800 1250 -1600 1650
rect -1550 1850 -1450 1900
rect -1550 1600 -1450 1650
rect -1400 1850 -1200 1900
rect -1400 1650 -1350 1850
rect -1250 1650 -1200 1850
rect -1800 1050 -1750 1250
rect -1650 1050 -1600 1250
rect -1800 1000 -1600 1050
rect -2850 850 -2800 950
rect -2500 850 -2150 950
rect -1850 850 -1800 950
rect -1750 750 -1600 1000
rect -2350 650 -2150 700
rect -2350 450 -2300 650
rect -2200 450 -2150 650
rect -2350 400 -2150 450
rect -1850 650 -1600 750
rect -1850 450 -1800 650
rect -1700 600 -1600 650
rect -1400 1250 -1200 1650
rect -1400 1050 -1350 1250
rect -1250 1050 -1200 1250
rect -1400 1000 -1200 1050
rect -800 1850 -600 1900
rect -800 1650 -750 1850
rect -650 1650 -600 1850
rect -800 1250 -600 1650
rect -800 1050 -750 1250
rect -650 1050 -600 1250
rect -800 1000 -600 1050
rect -150 1850 50 1950
rect -150 1650 -100 1850
rect 0 1650 50 1850
rect -150 1250 50 1650
rect 100 1850 200 1900
rect 100 1600 200 1650
rect -150 1050 -100 1250
rect 0 1050 50 1250
rect -150 1000 50 1050
rect -1400 750 -1250 1000
rect -1200 850 -1150 950
rect -850 850 -500 950
rect -200 850 -150 950
rect -1400 650 -1150 750
rect -1400 600 -1300 650
rect -1700 450 -1650 600
rect -1850 400 -1650 450
rect -1350 450 -1300 600
rect -1200 450 -1150 650
rect -1350 400 -1150 450
rect -850 650 -650 700
rect -850 450 -800 650
rect -700 450 -650 650
rect -850 400 -650 450
rect -2100 350 -900 400
rect -1900 250 -1100 350
rect -2100 200 -900 250
rect -1650 150 -1350 200
rect -1650 0 300 150
<< viali >>
rect -3000 6450 -2900 6650
rect -100 6450 0 6650
rect -1750 2850 -1650 3050
rect -1350 2850 -1250 3050
rect -2800 850 -2500 950
rect -2150 850 -1850 950
rect -2300 450 -2200 650
rect -1150 850 -850 950
rect -500 850 -200 950
rect -800 450 -700 650
<< metal1 >>
rect -3300 6650 300 6900
rect -3300 6450 -3000 6650
rect -2900 6450 -100 6650
rect 0 6450 300 6650
rect -3300 6100 300 6450
rect -1800 3050 -1200 3100
rect -1800 2850 -1750 3050
rect -1650 2850 -1350 3050
rect -1250 2850 -1200 3050
rect -1800 1000 -1200 2850
rect -3300 950 300 1000
rect -3300 850 -2800 950
rect -2500 850 -2150 950
rect -1850 850 -1150 950
rect -850 850 -500 950
rect -200 850 300 950
rect -3300 650 300 850
rect -3300 450 -2300 650
rect -2200 450 -800 650
rect -700 450 300 650
rect -3300 200 300 450
<< labels >>
rlabel locali 300 7000 300 7000 3 Vbp
port 1 e
rlabel metal1 300 6500 300 6500 3 VDD
port 2 e
rlabel locali 300 50 300 50 3 Vbn2
port 3 e
rlabel metal1 300 600 300 600 3 GND
port 4 e
<< end >>
