magic
tech sky130A
timestamp 1759703914
<< locali >>
rect 545 810 565 830
rect 915 810 935 830
rect 1285 810 1305 830
rect 1655 810 1675 830
rect -10 745 10 765
rect 1655 535 1675 555
<< metal1 >>
rect -10 460 10 770
rect -10 110 10 405
rect -10 -5 195 35
use d_ff  d_ff_0
timestamp 1759703914
transform 1 0 400 0 1 130
box -205 -135 165 700
use d_ff  d_ff_1
timestamp 1759703914
transform 1 0 770 0 1 130
box -205 -135 165 700
use d_ff  d_ff_2
timestamp 1759703914
transform 1 0 1140 0 1 130
box -205 -135 165 700
use d_ff  d_ff_3
timestamp 1759703914
transform 1 0 1510 0 1 130
box -205 -135 165 700
use inverter  inverter_0
timestamp 1759518789
transform 1 0 110 0 1 310
box -120 -200 100 520
<< labels >>
rlabel metal1 -10 15 -10 15 7 clk
port 0 w
rlabel locali -10 755 -10 755 7 D
port 1 w
rlabel locali 555 830 555 830 1 Q0
port 2 n
rlabel locali 925 830 925 830 1 Q1
port 3 n
rlabel locali 1295 830 1295 830 1 Q2
port 4 n
rlabel locali 1665 830 1665 830 1 Q3
port 5 n
rlabel metal1 -10 610 -10 610 7 VP
port 6 w
rlabel metal1 -10 255 -10 255 7 VN
port 7 w
rlabel locali 1675 545 1675 545 3 Qn3
port 8 e
<< end >>
