magic
tech sky130A
timestamp 1762058210
<< nwell >>
rect -2210 -270 -705 320
<< nmos >>
rect -2190 -845 -1890 -445
rect -1640 -845 -1340 -445
rect -1090 -845 -790 -445
rect 55 -815 1055 185
rect -5100 -1545 -4800 -1145
rect -4770 -1545 -4470 -1145
rect -4440 -1545 -4140 -1145
rect -4110 -1545 -3810 -1145
rect -3780 -1545 -3480 -1145
rect -3450 -1545 -3150 -1145
rect -3120 -1545 -2820 -1145
rect -2790 -1545 -2490 -1145
rect -2460 -1545 -2160 -1145
rect -2130 -1545 -1830 -1145
rect -1800 -1545 -1500 -1145
rect -1470 -1545 -1170 -1145
rect -1140 -1545 -840 -1145
rect -810 -1545 -510 -1145
rect -480 -1545 -180 -1145
rect -150 -1545 150 -1145
rect 180 -1545 480 -1145
rect 510 -1545 810 -1145
rect 840 -1545 1140 -1145
rect 1170 -1545 1470 -1145
<< pmos >>
rect -2190 -200 -1890 200
rect -1825 -200 -1525 200
rect -1365 -200 -1065 200
rect -1025 -200 -725 200
<< ndiff >>
rect 55 220 1055 235
rect 55 200 70 220
rect 1040 200 1055 220
rect 55 185 1055 200
rect -2190 -410 -1890 -395
rect -2190 -430 -2175 -410
rect -1905 -430 -1890 -410
rect -2190 -445 -1890 -430
rect -1640 -410 -1340 -395
rect -1640 -430 -1625 -410
rect -1355 -430 -1340 -410
rect -1640 -445 -1340 -430
rect -1090 -410 -790 -395
rect -1090 -430 -1075 -410
rect -805 -430 -790 -410
rect -1090 -445 -790 -430
rect 55 -830 1055 -815
rect -2190 -860 -1890 -845
rect -2190 -880 -2175 -860
rect -1905 -880 -1890 -860
rect -2190 -895 -1890 -880
rect -1640 -860 -1340 -845
rect -1640 -880 -1625 -860
rect -1355 -880 -1340 -860
rect -1640 -895 -1340 -880
rect -1090 -860 -790 -845
rect -1090 -880 -1075 -860
rect -805 -880 -790 -860
rect -1090 -885 -790 -880
rect 55 -850 70 -830
rect 1040 -850 1055 -830
rect 55 -865 1055 -850
rect -5100 -1110 -4800 -1095
rect -5100 -1130 -5085 -1110
rect -4815 -1130 -4800 -1110
rect -5100 -1145 -4800 -1130
rect -4770 -1110 -4470 -1095
rect -4770 -1130 -4755 -1110
rect -4485 -1130 -4470 -1110
rect -4770 -1145 -4470 -1130
rect -4440 -1110 -4140 -1095
rect -4440 -1130 -4425 -1110
rect -4155 -1130 -4140 -1110
rect -4440 -1145 -4140 -1130
rect -4110 -1110 -3810 -1095
rect -4110 -1130 -4095 -1110
rect -3825 -1130 -3810 -1110
rect -4110 -1145 -3810 -1130
rect -3780 -1110 -3480 -1095
rect -3780 -1130 -3765 -1110
rect -3495 -1130 -3480 -1110
rect -3780 -1145 -3480 -1130
rect -3450 -1110 -3150 -1095
rect -3450 -1130 -3435 -1110
rect -3165 -1130 -3150 -1110
rect -3450 -1145 -3150 -1130
rect -3120 -1110 -2820 -1095
rect -3120 -1130 -3105 -1110
rect -2835 -1130 -2820 -1110
rect -3120 -1145 -2820 -1130
rect -2790 -1110 -2490 -1095
rect -2790 -1130 -2775 -1110
rect -2505 -1130 -2490 -1110
rect -2790 -1145 -2490 -1130
rect -2460 -1110 -2160 -1095
rect -2460 -1130 -2445 -1110
rect -2175 -1130 -2160 -1110
rect -2460 -1145 -2160 -1130
rect -2130 -1110 -1830 -1095
rect -2130 -1130 -2115 -1110
rect -1845 -1130 -1830 -1110
rect -2130 -1145 -1830 -1130
rect -1800 -1110 -1500 -1095
rect -1800 -1130 -1785 -1110
rect -1515 -1130 -1500 -1110
rect -1800 -1145 -1500 -1130
rect -1470 -1110 -1170 -1095
rect -1470 -1130 -1455 -1110
rect -1185 -1130 -1170 -1110
rect -1470 -1145 -1170 -1130
rect -1140 -1110 -840 -1095
rect -1140 -1130 -1125 -1110
rect -855 -1130 -840 -1110
rect -1140 -1145 -840 -1130
rect -810 -1110 -510 -1095
rect -810 -1130 -795 -1110
rect -525 -1130 -510 -1110
rect -810 -1145 -510 -1130
rect -480 -1110 -180 -1095
rect -480 -1130 -465 -1110
rect -195 -1130 -180 -1110
rect -480 -1145 -180 -1130
rect -150 -1110 150 -1095
rect -150 -1130 -135 -1110
rect 135 -1130 150 -1110
rect -150 -1145 150 -1130
rect 180 -1110 480 -1095
rect 180 -1130 195 -1110
rect 465 -1130 480 -1110
rect 180 -1145 480 -1130
rect 510 -1110 810 -1095
rect 510 -1130 525 -1110
rect 795 -1130 810 -1110
rect 510 -1145 810 -1130
rect 840 -1110 1140 -1095
rect 840 -1130 855 -1110
rect 1125 -1130 1140 -1110
rect 840 -1145 1140 -1130
rect 1170 -1110 1470 -1095
rect 1170 -1130 1185 -1110
rect 1455 -1130 1470 -1110
rect 1170 -1145 1470 -1130
rect -5100 -1560 -4800 -1545
rect -5100 -1580 -5085 -1560
rect -4815 -1580 -4800 -1560
rect -5100 -1595 -4800 -1580
rect -4770 -1560 -4470 -1545
rect -4770 -1580 -4755 -1560
rect -4485 -1580 -4470 -1560
rect -4770 -1595 -4470 -1580
rect -4440 -1560 -4140 -1545
rect -4440 -1580 -4425 -1560
rect -4155 -1580 -4140 -1560
rect -4440 -1595 -4140 -1580
rect -4110 -1560 -3810 -1545
rect -4110 -1580 -4095 -1560
rect -3825 -1580 -3810 -1560
rect -4110 -1595 -3810 -1580
rect -3780 -1560 -3480 -1545
rect -3780 -1580 -3765 -1560
rect -3495 -1580 -3480 -1560
rect -3780 -1595 -3480 -1580
rect -3450 -1560 -3150 -1545
rect -3450 -1580 -3435 -1560
rect -3165 -1580 -3150 -1560
rect -3450 -1595 -3150 -1580
rect -3120 -1560 -2820 -1545
rect -3120 -1580 -3105 -1560
rect -2835 -1580 -2820 -1560
rect -3120 -1595 -2820 -1580
rect -2790 -1560 -2490 -1545
rect -2790 -1580 -2775 -1560
rect -2505 -1580 -2490 -1560
rect -2790 -1595 -2490 -1580
rect -2460 -1560 -2160 -1545
rect -2460 -1580 -2445 -1560
rect -2175 -1580 -2160 -1560
rect -2460 -1595 -2160 -1580
rect -2130 -1560 -1830 -1545
rect -2130 -1580 -2115 -1560
rect -1845 -1580 -1830 -1560
rect -2130 -1595 -1830 -1580
rect -1800 -1560 -1500 -1545
rect -1800 -1580 -1785 -1560
rect -1515 -1580 -1500 -1560
rect -1800 -1595 -1500 -1580
rect -1470 -1560 -1170 -1545
rect -1470 -1580 -1455 -1560
rect -1185 -1580 -1170 -1560
rect -1470 -1595 -1170 -1580
rect -1140 -1560 -840 -1545
rect -1140 -1580 -1125 -1560
rect -855 -1580 -840 -1560
rect -1140 -1595 -840 -1580
rect -810 -1560 -510 -1545
rect -810 -1580 -795 -1560
rect -525 -1580 -510 -1560
rect -810 -1595 -510 -1580
rect -480 -1560 -180 -1545
rect -480 -1580 -465 -1560
rect -195 -1580 -180 -1560
rect -480 -1595 -180 -1580
rect -150 -1560 150 -1545
rect -150 -1580 -135 -1560
rect 135 -1580 150 -1560
rect -150 -1595 150 -1580
rect 180 -1560 480 -1545
rect 180 -1580 195 -1560
rect 465 -1580 480 -1560
rect 180 -1595 480 -1580
rect 510 -1560 810 -1545
rect 510 -1580 525 -1560
rect 795 -1580 810 -1560
rect 510 -1595 810 -1580
rect 840 -1560 1140 -1545
rect 840 -1580 855 -1560
rect 1125 -1580 1140 -1560
rect 840 -1595 1140 -1580
rect 1170 -1560 1470 -1545
rect 1170 -1580 1185 -1560
rect 1455 -1580 1470 -1560
rect 1170 -1595 1470 -1580
<< pdiff >>
rect -2190 235 -1890 250
rect -2190 215 -2175 235
rect -1905 215 -1890 235
rect -2190 200 -1890 215
rect -1825 235 -1525 250
rect -1825 215 -1810 235
rect -1540 215 -1525 235
rect -1825 200 -1525 215
rect -1365 235 -1065 250
rect -1365 215 -1350 235
rect -1080 215 -1065 235
rect -1365 200 -1065 215
rect -1025 235 -725 250
rect -1025 215 -1010 235
rect -740 215 -725 235
rect -1025 200 -725 215
rect -2190 -215 -1890 -200
rect -2190 -235 -2170 -215
rect -1905 -235 -1890 -215
rect -2190 -250 -1890 -235
rect -1825 -215 -1525 -200
rect -1825 -235 -1805 -215
rect -1540 -235 -1525 -215
rect -1825 -250 -1525 -235
rect -1365 -215 -1065 -200
rect -1365 -235 -1345 -215
rect -1080 -235 -1065 -215
rect -1365 -250 -1065 -235
rect -1025 -215 -725 -200
rect -1025 -235 -1005 -215
rect -740 -235 -725 -215
rect -1025 -250 -725 -235
<< ndiffc >>
rect 70 200 1040 220
rect -2175 -430 -1905 -410
rect -1625 -430 -1355 -410
rect -1075 -430 -805 -410
rect -2175 -880 -1905 -860
rect -1625 -880 -1355 -860
rect -1075 -880 -805 -860
rect 70 -850 1040 -830
rect -5085 -1130 -4815 -1110
rect -4755 -1130 -4485 -1110
rect -4425 -1130 -4155 -1110
rect -4095 -1130 -3825 -1110
rect -3765 -1130 -3495 -1110
rect -3435 -1130 -3165 -1110
rect -3105 -1130 -2835 -1110
rect -2775 -1130 -2505 -1110
rect -2445 -1130 -2175 -1110
rect -2115 -1130 -1845 -1110
rect -1785 -1130 -1515 -1110
rect -1455 -1130 -1185 -1110
rect -1125 -1130 -855 -1110
rect -795 -1130 -525 -1110
rect -465 -1130 -195 -1110
rect -135 -1130 135 -1110
rect 195 -1130 465 -1110
rect 525 -1130 795 -1110
rect 855 -1130 1125 -1110
rect 1185 -1130 1455 -1110
rect -5085 -1580 -4815 -1560
rect -4755 -1580 -4485 -1560
rect -4425 -1580 -4155 -1560
rect -4095 -1580 -3825 -1560
rect -3765 -1580 -3495 -1560
rect -3435 -1580 -3165 -1560
rect -3105 -1580 -2835 -1560
rect -2775 -1580 -2505 -1560
rect -2445 -1580 -2175 -1560
rect -2115 -1580 -1845 -1560
rect -1785 -1580 -1515 -1560
rect -1455 -1580 -1185 -1560
rect -1125 -1580 -855 -1560
rect -795 -1580 -525 -1560
rect -465 -1580 -195 -1560
rect -135 -1580 135 -1560
rect 195 -1580 465 -1560
rect 525 -1580 795 -1560
rect 855 -1580 1125 -1560
rect 1185 -1580 1455 -1560
<< pdiffc >>
rect -2175 215 -1905 235
rect -1810 215 -1540 235
rect -1350 215 -1080 235
rect -1010 215 -740 235
rect -2170 -235 -1905 -215
rect -1805 -235 -1540 -215
rect -1345 -235 -1080 -215
rect -1005 -235 -740 -215
<< psubdiff >>
rect 55 270 1055 285
rect 55 250 70 270
rect 1040 250 1055 270
rect 55 235 1055 250
rect -2190 -910 -1890 -895
rect -2190 -930 -2175 -910
rect -1905 -930 -1890 -910
rect -2190 -945 -1890 -930
rect -1640 -910 -1340 -895
rect -1640 -930 -1625 -910
rect -1355 -930 -1340 -910
rect -1640 -945 -1340 -930
rect -1090 -900 -790 -885
rect -1090 -920 -1075 -900
rect -805 -920 -790 -900
rect 55 -880 1055 -865
rect 55 -900 70 -880
rect 1040 -900 1055 -880
rect 55 -915 1055 -900
rect -1090 -935 -790 -920
rect -4110 -1665 -3810 -1650
rect -4110 -1685 -4095 -1665
rect -3830 -1685 -3810 -1665
rect -4110 -1700 -3810 -1685
rect -300 -1665 0 -1650
rect -300 -1685 -285 -1665
rect -20 -1685 0 -1665
rect -300 -1700 0 -1685
rect -1831 -1770 -1611 -1755
rect -1831 -1790 -1816 -1770
rect -1631 -1790 -1611 -1770
rect -1831 -1805 -1611 -1790
<< nsubdiff >>
rect -2190 285 -1890 300
rect -2190 265 -2175 285
rect -1900 265 -1890 285
rect -2190 250 -1890 265
rect -1825 285 -1525 300
rect -1825 265 -1810 285
rect -1535 265 -1525 285
rect -1825 250 -1525 265
rect -1365 285 -1065 300
rect -1365 265 -1350 285
rect -1075 265 -1065 285
rect -1365 250 -1065 265
rect -1025 285 -725 300
rect -1025 265 -1010 285
rect -735 265 -725 285
rect -1025 250 -725 265
<< psubdiffcont >>
rect 70 250 1040 270
rect -2175 -930 -1905 -910
rect -1625 -930 -1355 -910
rect -1075 -920 -805 -900
rect 70 -900 1040 -880
rect -4095 -1685 -3830 -1665
rect -285 -1685 -20 -1665
rect -1816 -1790 -1631 -1770
<< nsubdiffcont >>
rect -2175 265 -1900 285
rect -1810 265 -1535 285
rect -1350 265 -1075 285
rect -1010 265 -735 285
<< poly >>
rect -2205 -175 -2190 200
rect -2235 -200 -2190 -175
rect -1890 -200 -1825 200
rect -1525 -200 -1510 200
rect -1380 -175 -1365 200
rect -1455 -200 -1365 -175
rect -1065 -200 -1025 200
rect -725 -140 -710 200
rect 40 -140 55 185
rect -725 -150 55 -140
rect -725 -190 -700 -150
rect -660 -190 55 -150
rect -725 -200 55 -190
rect -2235 -285 -2210 -200
rect -1455 -265 -1430 -200
rect -2185 -275 -2140 -265
rect -2185 -285 -2175 -275
rect -2235 -300 -2175 -285
rect -2150 -300 -2140 -275
rect -2235 -310 -2140 -300
rect -1575 -275 -1430 -265
rect -1575 -300 -1565 -275
rect -1540 -290 -1430 -275
rect -1540 -300 -1530 -290
rect -1575 -310 -1530 -300
rect -775 -410 -735 -400
rect -775 -430 -765 -410
rect -745 -430 -735 -410
rect -775 -445 -735 -430
rect -2220 -820 -2190 -445
rect -2425 -845 -2190 -820
rect -1890 -845 -1860 -445
rect -1670 -845 -1640 -445
rect -1340 -845 -1090 -445
rect -790 -455 -735 -445
rect -790 -845 -760 -455
rect 40 -815 55 -200
rect 1055 -815 1070 185
rect -2425 -1020 -2400 -845
rect -2460 -1030 -2400 -1020
rect -2460 -1070 -2450 -1030
rect -2425 -1050 -2400 -1030
rect -2410 -1070 -2400 -1050
rect -2460 -1080 -2400 -1070
rect -5115 -1545 -5100 -1145
rect -4800 -1545 -4770 -1145
rect -4470 -1545 -4440 -1145
rect -4140 -1545 -4110 -1145
rect -3810 -1545 -3780 -1145
rect -3480 -1545 -3450 -1145
rect -3150 -1545 -3120 -1145
rect -2820 -1545 -2790 -1145
rect -2490 -1545 -2460 -1145
rect -2160 -1545 -2130 -1145
rect -1830 -1545 -1800 -1145
rect -1500 -1545 -1470 -1145
rect -1170 -1545 -1140 -1145
rect -840 -1545 -810 -1145
rect -510 -1545 -480 -1145
rect -180 -1545 -150 -1145
rect 150 -1545 180 -1145
rect 480 -1545 510 -1145
rect 810 -1545 840 -1145
rect 1140 -1545 1170 -1145
rect 1470 -1155 1545 -1145
rect 1470 -1195 1495 -1155
rect 1535 -1195 1545 -1155
rect 1470 -1205 1545 -1195
rect 1470 -1545 1485 -1205
<< polycont >>
rect -700 -190 -660 -150
rect -2175 -300 -2150 -275
rect -1565 -300 -1540 -275
rect -765 -430 -745 -410
rect -2450 -1050 -2425 -1030
rect -2450 -1070 -2410 -1050
rect 1495 -1195 1535 -1155
<< xpolycontact >>
rect -3785 -1890 -3565 -1855
rect -1831 -1890 -1611 -1855
<< ppolyres >>
rect -3565 -1890 -1831 -1855
<< locali >>
rect -2190 285 -1890 300
rect -2190 265 -2175 285
rect -1900 265 -1890 285
rect -2190 235 -1890 265
rect -2190 215 -2175 235
rect -1905 215 -1890 235
rect -2190 200 -1890 215
rect -1825 285 -1525 300
rect -1825 265 -1810 285
rect -1535 265 -1525 285
rect -1825 235 -1525 265
rect -1825 215 -1810 235
rect -1540 215 -1525 235
rect -1825 200 -1525 215
rect -1365 285 -1065 300
rect -1365 265 -1350 285
rect -1075 265 -1065 285
rect -1365 235 -1065 265
rect -1365 215 -1350 235
rect -1080 215 -1065 235
rect -1365 200 -1065 215
rect -1025 285 -725 300
rect -1025 265 -1010 285
rect -735 265 -725 285
rect -1025 235 -725 265
rect -1025 215 -1010 235
rect -740 215 -725 235
rect -1025 200 -725 215
rect -650 -140 -630 325
rect -710 -150 -630 -140
rect -710 -190 -700 -150
rect -660 -190 -630 -150
rect -710 -200 -630 -190
rect -2185 -215 -1895 -205
rect -2185 -235 -2170 -215
rect -1905 -235 -1895 -215
rect -2185 -245 -1895 -235
rect -1820 -215 -1530 -205
rect -1820 -235 -1805 -215
rect -1540 -235 -1530 -215
rect -1820 -245 -1530 -235
rect -1360 -215 -1070 -205
rect -1360 -235 -1345 -215
rect -1080 -235 -1070 -215
rect -1360 -245 -1070 -235
rect -1020 -215 -730 -205
rect -1020 -235 -1005 -215
rect -740 -235 -730 -215
rect -1020 -245 -730 -235
rect -2185 -275 -2140 -245
rect -2185 -300 -2175 -275
rect -2150 -300 -2140 -275
rect -2185 -400 -2140 -300
rect -1575 -275 -1530 -245
rect -1575 -300 -1565 -275
rect -1540 -300 -1530 -275
rect -1575 -400 -1530 -300
rect -2220 -410 -1860 -400
rect -2220 -430 -2175 -410
rect -1905 -430 -1860 -410
rect -2220 -440 -1860 -430
rect -1670 -410 -1310 -400
rect -1670 -430 -1625 -410
rect -1355 -430 -1310 -410
rect -1670 -440 -1310 -430
rect -2220 -860 -1860 -850
rect -2220 -880 -2175 -860
rect -1905 -880 -1860 -860
rect -2220 -890 -1860 -880
rect -1670 -860 -1310 -850
rect -1670 -880 -1625 -860
rect -1355 -880 -1310 -860
rect -1670 -890 -1310 -880
rect -2190 -910 -1890 -890
rect -2190 -930 -2175 -910
rect -1905 -930 -1890 -910
rect -2190 -945 -1890 -930
rect -1640 -910 -1340 -890
rect -1640 -930 -1625 -910
rect -1355 -930 -1340 -910
rect -1640 -945 -1340 -930
rect -2460 -1030 -2400 -1020
rect -2460 -1070 -2450 -1030
rect -2425 -1050 -2400 -1030
rect -2410 -1070 -2400 -1050
rect -2460 -1080 -2400 -1070
rect -2460 -1100 -2440 -1080
rect -1230 -1100 -1190 -245
rect -1020 -400 -980 -245
rect -565 -400 -545 325
rect 60 270 1050 280
rect 60 250 70 270
rect 1040 250 1050 270
rect 60 220 1050 250
rect 60 200 70 220
rect 1040 200 1050 220
rect 60 190 1050 200
rect -1120 -410 -545 -400
rect -1120 -430 -1075 -410
rect -805 -430 -765 -410
rect -745 -420 -545 -410
rect -745 -430 -735 -420
rect -1120 -440 -735 -430
rect 60 -830 1050 -820
rect 60 -850 70 -830
rect 1040 -850 1050 -830
rect -1120 -860 -760 -850
rect -1120 -880 -1075 -860
rect -805 -880 -760 -860
rect -1120 -890 -760 -880
rect 60 -880 1050 -850
rect -1090 -900 -790 -890
rect -1090 -920 -1075 -900
rect -805 -920 -790 -900
rect 60 -900 70 -880
rect 1040 -900 1050 -880
rect 60 -910 1050 -900
rect -1090 -935 -790 -920
rect -5095 -1110 1545 -1100
rect -5095 -1130 -5085 -1110
rect -4815 -1130 -4755 -1110
rect -4485 -1130 -4425 -1110
rect -4155 -1130 -4095 -1110
rect -3825 -1130 -3765 -1110
rect -3495 -1130 -3435 -1110
rect -3165 -1130 -3105 -1110
rect -2835 -1130 -2775 -1110
rect -2505 -1130 -2445 -1110
rect -2175 -1130 -2115 -1110
rect -1845 -1130 -1785 -1110
rect -1515 -1130 -1455 -1110
rect -1185 -1130 -1125 -1110
rect -855 -1130 -795 -1110
rect -525 -1130 -465 -1110
rect -195 -1130 -135 -1110
rect 135 -1130 195 -1110
rect 465 -1130 525 -1110
rect 795 -1130 855 -1110
rect 1125 -1130 1185 -1110
rect 1455 -1130 1545 -1110
rect -5095 -1140 1545 -1130
rect 1485 -1155 1545 -1140
rect 1485 -1195 1495 -1155
rect 1535 -1195 1545 -1155
rect 1485 -1205 1545 -1195
rect -5095 -1560 1465 -1550
rect -5095 -1580 -5085 -1560
rect -4815 -1580 -4755 -1560
rect -4485 -1580 -4425 -1560
rect -4155 -1580 -4095 -1560
rect -3825 -1580 -3765 -1560
rect -3495 -1580 -3435 -1560
rect -3165 -1580 -3105 -1560
rect -2835 -1580 -2775 -1560
rect -2505 -1580 -2445 -1560
rect -2175 -1580 -2115 -1560
rect -1845 -1580 -1785 -1560
rect -1515 -1580 -1455 -1560
rect -1185 -1580 -1125 -1560
rect -855 -1580 -795 -1560
rect -525 -1580 -465 -1560
rect -195 -1580 -135 -1560
rect 135 -1580 195 -1560
rect 465 -1580 525 -1560
rect 795 -1580 855 -1560
rect 1125 -1580 1185 -1560
rect 1455 -1580 1465 -1560
rect -5095 -1590 1465 -1580
rect -4105 -1665 -3815 -1655
rect -4105 -1685 -4095 -1665
rect -3830 -1685 -3815 -1665
rect -4105 -1695 -3815 -1685
rect -3785 -1855 -3565 -1590
rect -295 -1665 -5 -1655
rect -295 -1685 -285 -1665
rect -20 -1685 -5 -1665
rect -295 -1695 -5 -1685
rect -1826 -1770 -1616 -1760
rect -1826 -1790 -1816 -1770
rect -1631 -1790 -1616 -1770
rect -1826 -1855 -1616 -1790
<< viali >>
rect -2175 265 -1900 285
rect -1810 265 -1540 285
rect -1350 265 -1080 285
rect -1010 265 -740 285
rect -2175 -930 -1905 -910
rect -1625 -930 -1355 -910
rect 70 250 1040 270
rect -1075 -920 -805 -900
rect 70 -900 1040 -880
rect -4095 -1685 -3830 -1665
rect -285 -1685 -20 -1665
<< metal1 >>
rect -5115 285 -705 320
rect -5115 265 -2175 285
rect -1900 265 -1810 285
rect -1540 265 -1350 285
rect -1080 265 -1010 285
rect -740 265 -705 285
rect -5115 -715 -705 265
rect -165 270 1210 355
rect -165 250 70 270
rect 1040 250 1210 270
rect -2270 -900 -715 -785
rect -2270 -905 -1075 -900
rect -5115 -910 -1075 -905
rect -5115 -930 -2175 -910
rect -1905 -930 -1625 -910
rect -1355 -920 -1075 -910
rect -805 -905 -715 -900
rect -165 -880 1210 250
rect -165 -900 70 -880
rect 1040 -900 1210 -880
rect -165 -905 1210 -900
rect -805 -920 1585 -905
rect -1355 -930 1585 -920
rect -5115 -1665 1585 -930
rect -5115 -1685 -4095 -1665
rect -3830 -1685 -285 -1665
rect -20 -1685 1585 -1665
rect -5115 -1910 1585 -1685
<< labels >>
rlabel metal1 -5115 -965 -5115 -965 7 GND
port 3 w
rlabel metal1 -5115 -175 -5115 -175 7 VDD
port 2 w
rlabel locali -640 325 -640 325 1 Vbp
port 1 n
rlabel locali -555 325 -555 325 1 Vbn
port 0 n
<< properties >>
string MASKHINTS_RPM -3805 -1950 -1575 -1780
string MASKHINTS_URPM -3880 -2010 -1522 -1689
<< end >>
