magic
tech sky130A
timestamp 1762122866
<< nmos >>
rect 2800 7200 3000 8100
rect -200 6850 200 7150
rect 400 6850 800 7150
rect 900 7000 1300 7100
rect 1850 6250 2050 7150
rect 2300 6250 2500 7150
rect 2800 6250 3000 7150
rect -200 5900 200 6200
rect 400 5900 800 6200
rect 900 6050 1300 6150
rect 1850 5300 2050 6200
rect 2300 5300 2500 6200
rect 2800 5300 3000 6200
rect -200 4950 200 5250
rect 400 4950 800 5250
rect 900 5100 1300 5200
rect 1850 4350 2050 5250
rect 2300 4350 2500 5250
rect 2800 4350 3000 5250
rect -200 4000 200 4300
rect 400 4000 800 4300
rect 900 4150 1300 4250
rect 1850 3400 2050 4300
rect 2300 3400 2500 4300
rect 2800 3400 3000 4300
rect -200 3050 200 3350
rect 400 3050 800 3350
rect 900 3200 1300 3300
rect 1850 2450 2050 3350
rect 2300 2450 2500 3350
rect 2800 2450 3000 3350
rect -200 2100 200 2400
rect 400 2100 800 2400
rect 900 2250 1300 2350
rect 1850 1500 2050 2400
rect 2300 1500 2500 2400
rect 2800 1500 3000 2400
rect -200 1150 200 1450
rect 400 1150 800 1450
rect 900 1300 1300 1400
rect 2800 550 3000 1450
rect 2800 -400 3000 500
<< ndiff >>
rect 2550 8000 2800 8100
rect 2550 7300 2650 8000
rect 2700 7300 2800 8000
rect 2550 7200 2800 7300
rect 3000 8000 3250 8100
rect 3000 7300 3100 8000
rect 3150 7300 3250 8000
rect 3000 7200 3250 7300
rect -400 7050 -200 7150
rect -400 6950 -350 7050
rect -250 6950 -200 7050
rect -400 6850 -200 6950
rect 200 6850 400 7150
rect 800 7100 850 7150
rect 1600 7100 1850 7150
rect 800 7000 900 7100
rect 1300 7050 1850 7100
rect 1300 7000 1700 7050
rect 800 6850 850 7000
rect 1600 6800 1700 7000
rect 1650 6750 1700 6800
rect 1600 6350 1700 6750
rect 1750 6350 1850 7050
rect 1600 6250 1850 6350
rect 2050 6600 2300 7150
rect 2050 6300 2150 6600
rect 2200 6300 2300 6600
rect 2050 6250 2300 6300
rect 2500 7050 2800 7150
rect 2500 6350 2650 7050
rect 2700 6350 2800 7050
rect 2500 6250 2800 6350
rect 3000 7050 3250 7150
rect 3000 6350 3100 7050
rect 3150 6350 3250 7050
rect 3000 6250 3250 6350
rect -400 6100 -200 6200
rect -400 6000 -350 6100
rect -250 6000 -200 6100
rect -400 5900 -200 6000
rect 200 5900 400 6200
rect 800 6150 850 6200
rect 1600 6150 1850 6200
rect 800 6050 900 6150
rect 1300 6100 1850 6150
rect 1300 6050 1700 6100
rect 800 5900 850 6050
rect 1600 5850 1700 6050
rect 1650 5800 1700 5850
rect 1600 5400 1700 5800
rect 1750 5400 1850 6100
rect 1600 5300 1850 5400
rect 2050 5650 2300 6200
rect 2050 5350 2150 5650
rect 2200 5350 2300 5650
rect 2050 5300 2300 5350
rect 2500 6100 2800 6200
rect 2500 5400 2650 6100
rect 2700 5400 2800 6100
rect 2500 5300 2800 5400
rect 3000 6100 3250 6200
rect 3000 5400 3100 6100
rect 3150 5400 3250 6100
rect 3000 5300 3250 5400
rect -400 5150 -200 5250
rect -400 5050 -350 5150
rect -250 5050 -200 5150
rect -400 4950 -200 5050
rect 200 4950 400 5250
rect 800 5200 850 5250
rect 1600 5200 1850 5250
rect 800 5100 900 5200
rect 1300 5150 1850 5200
rect 1300 5100 1700 5150
rect 800 4950 850 5100
rect 1600 4900 1700 5100
rect 1650 4850 1700 4900
rect 1600 4450 1700 4850
rect 1750 4450 1850 5150
rect 1600 4350 1850 4450
rect 2050 4700 2300 5250
rect 2050 4400 2150 4700
rect 2200 4400 2300 4700
rect 2050 4350 2300 4400
rect 2500 5150 2800 5250
rect 2500 4450 2650 5150
rect 2700 4450 2800 5150
rect 2500 4350 2800 4450
rect 3000 5150 3250 5250
rect 3000 4450 3100 5150
rect 3150 4450 3250 5150
rect 3000 4350 3250 4450
rect -400 4200 -200 4300
rect -400 4100 -350 4200
rect -250 4100 -200 4200
rect -400 4000 -200 4100
rect 200 4000 400 4300
rect 800 4250 850 4300
rect 1600 4250 1850 4300
rect 800 4150 900 4250
rect 1300 4200 1850 4250
rect 1300 4150 1700 4200
rect 800 4000 850 4150
rect 1600 3950 1700 4150
rect 1650 3900 1700 3950
rect 1600 3500 1700 3900
rect 1750 3500 1850 4200
rect 1600 3400 1850 3500
rect 2050 3750 2300 4300
rect 2050 3450 2150 3750
rect 2200 3450 2300 3750
rect 2050 3400 2300 3450
rect 2500 4200 2800 4300
rect 2500 3500 2650 4200
rect 2700 3500 2800 4200
rect 2500 3400 2800 3500
rect 3000 4200 3250 4300
rect 3000 3500 3100 4200
rect 3150 3500 3250 4200
rect 3000 3400 3250 3500
rect -400 3250 -200 3350
rect -400 3150 -350 3250
rect -250 3150 -200 3250
rect -400 3050 -200 3150
rect 200 3050 400 3350
rect 800 3300 850 3350
rect 1600 3300 1850 3350
rect 800 3200 900 3300
rect 1300 3250 1850 3300
rect 1300 3200 1700 3250
rect 800 3050 850 3200
rect 1600 3000 1700 3200
rect 1650 2950 1700 3000
rect 1600 2550 1700 2950
rect 1750 2550 1850 3250
rect 1600 2450 1850 2550
rect 2050 2800 2300 3350
rect 2050 2500 2150 2800
rect 2200 2500 2300 2800
rect 2050 2450 2300 2500
rect 2500 3250 2800 3350
rect 2500 2550 2650 3250
rect 2700 2550 2800 3250
rect 2500 2450 2800 2550
rect 3000 3250 3250 3350
rect 3000 2550 3100 3250
rect 3150 2550 3250 3250
rect 3000 2450 3250 2550
rect -400 2300 -200 2400
rect -400 2200 -350 2300
rect -250 2200 -200 2300
rect -400 2100 -200 2200
rect 200 2100 400 2400
rect 800 2350 850 2400
rect 1600 2350 1850 2400
rect 800 2250 900 2350
rect 1300 2300 1850 2350
rect 1300 2250 1700 2300
rect 800 2100 850 2250
rect 1600 2050 1700 2250
rect 1650 2000 1700 2050
rect 1600 1600 1700 2000
rect 1750 1600 1850 2300
rect 1600 1500 1850 1600
rect 2050 1850 2300 2400
rect 2050 1550 2150 1850
rect 2200 1550 2300 1850
rect 2050 1500 2300 1550
rect 2500 2300 2800 2400
rect 2500 1600 2650 2300
rect 2700 1600 2800 2300
rect 2500 1500 2800 1600
rect 3000 2300 3250 2400
rect 3000 1600 3100 2300
rect 3150 1600 3250 2300
rect 3000 1500 3250 1600
rect -400 1350 -200 1450
rect -400 1250 -350 1350
rect -250 1250 -200 1350
rect -400 1150 -200 1250
rect 200 1150 400 1450
rect 800 1400 850 1450
rect 1600 1400 1800 1450
rect 800 1300 900 1400
rect 1300 1350 1800 1400
rect 1300 1300 1700 1350
rect 800 1150 850 1300
rect 1600 1100 1700 1300
rect 1650 1050 1700 1100
rect 1600 650 1700 1050
rect 1750 650 1800 1350
rect 2550 1350 2800 1450
rect 1600 550 1800 650
rect 2550 650 2650 1350
rect 2700 650 2800 1350
rect 2550 550 2800 650
rect 3000 1350 3250 1450
rect 3000 650 3100 1350
rect 3150 650 3250 1350
rect 3000 550 3250 650
rect 2550 400 2800 500
rect 2550 -300 2650 400
rect 2700 -300 2800 400
rect 2550 -400 2800 -300
rect 3000 400 3250 500
rect 3000 -300 3100 400
rect 3150 -300 3250 400
rect 3000 -400 3250 -300
<< ndiffc >>
rect 2650 7300 2700 8000
rect 3100 7300 3150 8000
rect -350 6950 -250 7050
rect 1700 6350 1750 7050
rect 2150 6300 2200 6600
rect 2650 6350 2700 7050
rect 3100 6350 3150 7050
rect -350 6000 -250 6100
rect 1700 5400 1750 6100
rect 2150 5350 2200 5650
rect 2650 5400 2700 6100
rect 3100 5400 3150 6100
rect -350 5050 -250 5150
rect 1700 4450 1750 5150
rect 2150 4400 2200 4700
rect 2650 4450 2700 5150
rect 3100 4450 3150 5150
rect -350 4100 -250 4200
rect 1700 3500 1750 4200
rect 2150 3450 2200 3750
rect 2650 3500 2700 4200
rect 3100 3500 3150 4200
rect -350 3150 -250 3250
rect 1700 2550 1750 3250
rect 2150 2500 2200 2800
rect 2650 2550 2700 3250
rect 3100 2550 3150 3250
rect -350 2200 -250 2300
rect 1700 1600 1750 2300
rect 2150 1550 2200 1850
rect 2650 1600 2700 2300
rect 3100 1600 3150 2300
rect -350 1250 -250 1350
rect 1700 650 1750 1350
rect 2650 650 2700 1350
rect 3100 650 3150 1350
rect 2650 -300 2700 400
rect 3100 -300 3150 400
<< psubdiff >>
rect 3250 8000 3500 8100
rect 3250 7300 3350 8000
rect 3400 7300 3500 8000
rect 3250 7200 3500 7300
rect -600 7050 -400 7150
rect -600 6950 -550 7050
rect -450 6950 -400 7050
rect -600 6850 -400 6950
rect 1350 6650 1600 6750
rect 1350 6350 1450 6650
rect 1500 6350 1600 6650
rect 1350 6250 1600 6350
rect -600 6100 -400 6200
rect -600 6000 -550 6100
rect -450 6000 -400 6100
rect -600 5900 -400 6000
rect 1350 5700 1600 5800
rect 1350 5400 1450 5700
rect 1500 5400 1600 5700
rect 1350 5300 1600 5400
rect 3250 6100 3500 6200
rect 3250 5400 3350 6100
rect 3400 5400 3500 6100
rect 3250 5300 3500 5400
rect -600 5150 -400 5250
rect -600 5050 -550 5150
rect -450 5050 -400 5150
rect -600 4950 -400 5050
rect 1350 4750 1600 4850
rect 1350 4450 1450 4750
rect 1500 4450 1600 4750
rect 1350 4350 1600 4450
rect -600 4200 -400 4300
rect -600 4100 -550 4200
rect -450 4100 -400 4200
rect -600 4000 -400 4100
rect 1350 3800 1600 3900
rect 1350 3500 1450 3800
rect 1500 3500 1600 3800
rect 1350 3400 1600 3500
rect 3250 4200 3500 4300
rect 3250 3500 3350 4200
rect 3400 3500 3500 4200
rect 3250 3400 3500 3500
rect -600 3250 -400 3350
rect -600 3150 -550 3250
rect -450 3150 -400 3250
rect -600 3050 -400 3150
rect 1350 2850 1600 2950
rect 1350 2550 1450 2850
rect 1500 2550 1600 2850
rect 1350 2450 1600 2550
rect -600 2300 -400 2400
rect -600 2200 -550 2300
rect -450 2200 -400 2300
rect -600 2100 -400 2200
rect 1350 1900 1600 2000
rect 1350 1600 1450 1900
rect 1500 1600 1600 1900
rect 1350 1500 1600 1600
rect 3250 2300 3500 2400
rect 3250 1600 3350 2300
rect 3400 1600 3500 2300
rect 3250 1500 3500 1600
rect -600 1350 -400 1450
rect -600 1250 -550 1350
rect -450 1250 -400 1350
rect -600 1150 -400 1250
rect 1350 950 1600 1050
rect 1350 650 1450 950
rect 1500 650 1600 950
rect 1350 550 1600 650
rect 3250 400 3500 500
rect 3250 -300 3350 400
rect 3400 -300 3500 400
rect 3250 -400 3500 -300
<< psubdiffcont >>
rect 3350 7300 3400 8000
rect -550 6950 -450 7050
rect 1450 6350 1500 6650
rect -550 6000 -450 6100
rect 1450 5400 1500 5700
rect 3350 5400 3400 6100
rect -550 5050 -450 5150
rect 1450 4450 1500 4750
rect -550 4100 -450 4200
rect 1450 3500 1500 3800
rect 3350 3500 3400 4200
rect -550 3150 -450 3250
rect 1450 2550 1500 2850
rect -550 2200 -450 2300
rect 1450 1600 1500 1900
rect 3350 1600 3400 2300
rect -550 1250 -450 1350
rect 1450 650 1500 950
rect 3350 -300 3400 400
<< poly >>
rect 1850 8300 2050 8350
rect -200 8250 200 8300
rect -200 8150 -150 8250
rect 150 8150 200 8250
rect -200 7150 200 8150
rect 400 8250 800 8300
rect 400 8150 450 8250
rect 750 8150 800 8250
rect 400 7150 800 8150
rect 1850 8200 1900 8300
rect 2000 8200 2050 8300
rect 1850 7150 2050 8200
rect 2300 8300 2500 8350
rect 2300 8200 2350 8300
rect 2450 8200 2500 8300
rect 2300 7150 2500 8200
rect 2800 8300 3000 8350
rect 2800 8200 2850 8300
rect 2950 8200 3000 8300
rect 2800 8100 3000 8200
rect 2800 7150 3000 7200
rect 900 7100 1300 7150
rect -200 6200 200 6850
rect 400 6200 800 6850
rect 900 6400 1300 7000
rect 900 6300 950 6400
rect 1250 6300 1300 6400
rect 900 6250 1300 6300
rect 1850 6200 2050 6250
rect 2300 6200 2500 6250
rect 2800 6200 3000 6250
rect 900 6150 1300 6200
rect -200 5250 200 5900
rect 400 5250 800 5900
rect 900 5450 1300 6050
rect 900 5350 950 5450
rect 1250 5350 1300 5450
rect 900 5300 1300 5350
rect 1850 5250 2050 5300
rect 2300 5250 2500 5300
rect 2800 5250 3000 5300
rect 900 5200 1300 5250
rect -200 4300 200 4950
rect 400 4300 800 4950
rect 900 4500 1300 5100
rect 900 4400 950 4500
rect 1250 4400 1300 4500
rect 900 4350 1300 4400
rect 1850 4300 2050 4350
rect 2300 4300 2500 4350
rect 2800 4300 3000 4350
rect 900 4250 1300 4300
rect -200 3350 200 4000
rect 400 3350 800 4000
rect 900 3550 1300 4150
rect 900 3450 950 3550
rect 1250 3450 1300 3550
rect 900 3400 1300 3450
rect 1850 3350 2050 3400
rect 2300 3350 2500 3400
rect 2800 3350 3000 3400
rect 900 3300 1300 3350
rect -200 2400 200 3050
rect 400 2400 800 3050
rect 900 2600 1300 3200
rect 900 2500 950 2600
rect 1250 2500 1300 2600
rect 900 2450 1300 2500
rect 1850 2400 2050 2450
rect 2300 2400 2500 2450
rect 2800 2400 3000 2450
rect 900 2350 1300 2400
rect -200 1450 200 2100
rect 400 1450 800 2100
rect 900 1650 1300 2250
rect 900 1550 950 1650
rect 1250 1550 1300 1650
rect 900 1500 1300 1550
rect 900 1400 1300 1450
rect -200 1100 200 1150
rect 400 1100 800 1150
rect 900 700 1300 1300
rect 900 600 950 700
rect 1250 600 1300 700
rect 900 550 1300 600
rect 1850 950 2050 1500
rect 2300 950 2500 1500
rect 2800 1450 3000 1500
rect 2800 500 3000 550
rect 2800 -550 3000 -400
<< polycont >>
rect -150 8150 150 8250
rect 450 8150 750 8250
rect 1900 8200 2000 8300
rect 2350 8200 2450 8300
rect 2850 8200 2950 8300
rect 950 6300 1250 6400
rect 950 5350 1250 5450
rect 950 4400 1250 4500
rect 950 3450 1250 3550
rect 950 2500 1250 2600
rect 950 1550 1250 1650
rect 950 600 1250 700
<< locali >>
rect -650 8700 1850 8850
rect -650 8500 800 8650
rect -650 8300 200 8450
rect -200 8250 200 8300
rect -200 8150 -150 8250
rect 150 8150 200 8250
rect -200 8100 200 8150
rect 400 8250 800 8500
rect 400 8150 450 8250
rect 750 8150 800 8250
rect 1650 8350 1850 8700
rect 1650 8300 3000 8350
rect 1650 8200 1900 8300
rect 2000 8200 2350 8300
rect 2450 8200 2850 8300
rect 2950 8200 3000 8300
rect 1650 8150 3000 8200
rect 400 8100 800 8150
rect 2600 8000 2750 8050
rect 2600 7300 2650 8000
rect 2700 7300 2750 8000
rect 2600 7100 2750 7300
rect -550 7050 -250 7100
rect -450 6950 -350 7050
rect -550 6900 -250 6950
rect -400 6850 -250 6900
rect 1650 7050 2750 7100
rect 1650 6700 1700 7050
rect 1400 6650 1550 6700
rect -650 6400 1300 6450
rect -650 6300 950 6400
rect 1250 6300 1300 6400
rect 1400 6350 1450 6650
rect 1500 6350 1550 6650
rect 1400 6300 1550 6350
rect 1600 6350 1700 6700
rect 1750 6700 2650 7050
rect 1750 6350 1800 6700
rect 1600 6300 1800 6350
rect 2100 6600 2250 6650
rect 2100 6300 2150 6600
rect 2200 6300 2250 6600
rect 2600 6350 2650 6700
rect 2700 6350 2750 7050
rect 2600 6300 2750 6350
rect 3050 8000 3250 8050
rect 3050 7300 3100 8000
rect 3150 7300 3250 8000
rect 3050 7250 3250 7300
rect 3300 8000 3450 8050
rect 3300 7300 3350 8000
rect 3400 7300 3450 8000
rect 3300 7250 3450 7300
rect 3050 7050 3200 7250
rect 3050 6350 3100 7050
rect 3150 6350 3200 7050
rect -650 6250 1300 6300
rect -400 6150 -250 6200
rect 2100 6150 2250 6300
rect 3050 6150 3200 6350
rect -550 6100 -250 6150
rect -450 6000 -350 6100
rect -550 5950 -250 6000
rect -400 5900 -250 5950
rect 1650 6100 2750 6150
rect 1400 5700 1550 5750
rect -650 5450 1300 5500
rect -650 5350 950 5450
rect 1250 5350 1300 5450
rect 1400 5400 1450 5700
rect 1500 5400 1550 5700
rect 1400 5350 1550 5400
rect 1650 5400 1700 6100
rect 1750 5750 2650 6100
rect 1750 5400 1800 5750
rect 1650 5350 1800 5400
rect 2100 5650 2250 5700
rect 2100 5350 2150 5650
rect 2200 5350 2250 5650
rect 2600 5400 2650 5750
rect 2700 5400 2750 6100
rect 2600 5350 2750 5400
rect 3050 6100 3250 6150
rect 3050 5400 3100 6100
rect 3150 5400 3250 6100
rect 3050 5350 3250 5400
rect 3300 6100 3450 6150
rect 3300 5400 3350 6100
rect 3400 5400 3450 6100
rect 3300 5350 3450 5400
rect -650 5300 1300 5350
rect -400 5200 -250 5250
rect 2100 5200 2250 5350
rect -550 5150 -250 5200
rect -450 5050 -350 5150
rect -550 5000 -250 5050
rect -400 4950 -250 5000
rect 1650 5150 2750 5200
rect 1400 4750 1550 4800
rect -650 4500 1300 4550
rect -650 4400 950 4500
rect 1250 4400 1300 4500
rect 1400 4450 1450 4750
rect 1500 4450 1550 4750
rect 1400 4400 1550 4450
rect 1650 4450 1700 5150
rect 1750 4800 2650 5150
rect 1750 4450 1800 4800
rect 1650 4400 1800 4450
rect 2100 4700 2250 4750
rect 2100 4400 2150 4700
rect 2200 4400 2250 4700
rect 2600 4450 2650 4800
rect 2700 4450 2750 5150
rect 2600 4400 2750 4450
rect 3050 5150 3200 5350
rect 3050 4450 3100 5150
rect 3150 4450 3200 5150
rect -650 4350 1300 4400
rect -400 4250 -250 4300
rect 2100 4250 2250 4400
rect 3050 4250 3200 4450
rect -550 4200 -250 4250
rect -450 4100 -350 4200
rect -550 4050 -250 4100
rect -400 4000 -250 4050
rect 1650 4200 2750 4250
rect 1400 3800 1550 3850
rect -650 3550 1300 3600
rect -650 3450 950 3550
rect 1250 3450 1300 3550
rect 1400 3500 1450 3800
rect 1500 3500 1550 3800
rect 1400 3450 1550 3500
rect 1650 3500 1700 4200
rect 1750 3850 2650 4200
rect 1750 3500 1800 3850
rect 1650 3450 1800 3500
rect 2100 3750 2250 3800
rect 2100 3450 2150 3750
rect 2200 3450 2250 3750
rect 2600 3500 2650 3850
rect 2700 3500 2750 4200
rect 2600 3450 2750 3500
rect 3050 4200 3250 4250
rect 3050 3500 3100 4200
rect 3150 3500 3250 4200
rect 3050 3450 3250 3500
rect 3300 4200 3450 4250
rect 3300 3500 3350 4200
rect 3400 3500 3450 4200
rect 3300 3450 3450 3500
rect -650 3400 1300 3450
rect -400 3300 -250 3350
rect 2100 3300 2250 3450
rect -550 3250 -250 3300
rect -450 3150 -350 3250
rect -550 3100 -250 3150
rect -400 3050 -250 3100
rect 1650 3250 2750 3300
rect 1400 2850 1550 2900
rect -650 2600 1300 2650
rect -650 2500 950 2600
rect 1250 2500 1300 2600
rect 1400 2550 1450 2850
rect 1500 2550 1550 2850
rect 1400 2500 1550 2550
rect 1650 2550 1700 3250
rect 1750 2900 2650 3250
rect 1750 2550 1800 2900
rect 1650 2500 1800 2550
rect 2100 2800 2250 2850
rect 2100 2500 2150 2800
rect 2200 2500 2250 2800
rect 2600 2550 2650 2900
rect 2700 2550 2750 3250
rect 2600 2500 2750 2550
rect 3050 3250 3200 3450
rect 3050 2550 3100 3250
rect 3150 2550 3200 3250
rect -650 2450 1300 2500
rect -400 2350 -250 2400
rect 2100 2350 2250 2500
rect 3050 2350 3200 2550
rect -550 2300 -250 2350
rect -450 2200 -350 2300
rect -550 2150 -250 2200
rect -400 2100 -250 2150
rect 1650 2300 2750 2350
rect 1400 1900 1550 1950
rect -650 1650 1300 1700
rect -650 1550 950 1650
rect 1250 1550 1300 1650
rect 1400 1600 1450 1900
rect 1500 1600 1550 1900
rect 1400 1550 1550 1600
rect 1650 1600 1700 2300
rect 1750 1950 2650 2300
rect 1750 1600 1800 1950
rect 1650 1550 1800 1600
rect 2100 1850 2250 1900
rect 2100 1550 2150 1850
rect 2200 1550 2250 1850
rect 2600 1600 2650 1950
rect 2700 1600 2750 2300
rect 2600 1550 2750 1600
rect 3050 2300 3250 2350
rect 3050 1600 3100 2300
rect 3150 1600 3250 2300
rect 3050 1550 3250 1600
rect 3300 2300 3450 2350
rect 3300 1600 3350 2300
rect 3400 1600 3450 2300
rect 3300 1550 3450 1600
rect -650 1500 1300 1550
rect -400 1400 -250 1450
rect 2100 1400 2250 1550
rect -550 1350 -250 1400
rect -450 1250 -350 1350
rect -550 1200 -250 1250
rect 1650 1350 2750 1400
rect 1400 950 1550 1000
rect -650 700 1300 750
rect -650 600 950 700
rect 1250 600 1300 700
rect 1400 650 1450 950
rect 1500 650 1550 950
rect 1400 600 1550 650
rect 1650 650 1700 1350
rect 1750 1000 2650 1350
rect 1750 650 1800 1000
rect 1650 600 1800 650
rect 2600 650 2650 1000
rect 2700 650 2750 1350
rect -650 550 1300 600
rect 2600 400 2750 650
rect 2600 -300 2650 400
rect 2700 -300 2750 400
rect 2600 -350 2750 -300
rect 3050 1350 3200 1400
rect 3050 650 3100 1350
rect 3150 650 3200 1350
rect 3050 400 3200 650
rect 3050 -300 3100 400
rect 3150 -300 3200 400
rect 3050 -450 3200 -300
rect 3300 400 3450 450
rect 3300 -300 3350 400
rect 3400 -300 3450 400
rect 3300 -350 3450 -300
rect 3050 -600 3550 -450
<< viali >>
rect -350 6950 -250 7050
rect 3100 7300 3150 8000
rect 3100 6350 3150 7050
rect -350 6000 -250 6100
rect 3100 5400 3150 6100
rect -350 5050 -250 5150
rect 3100 4450 3150 5150
rect -350 4100 -250 4200
rect 3100 3500 3150 4200
rect -350 3150 -250 3250
rect 3100 2550 3150 3250
rect -350 2200 -250 2300
rect 3100 1600 3150 2300
rect -350 1250 -250 1350
<< metal1 >>
rect -650 8000 3500 8100
rect -650 7300 3100 8000
rect 3150 7300 3500 8000
rect -650 7200 3500 7300
rect -550 7050 -200 7100
rect -550 6950 -350 7050
rect -250 6950 -200 7050
rect -550 6100 -200 6950
rect -550 6000 -350 6100
rect -250 6000 -200 6100
rect -550 5150 -200 6000
rect -550 5050 -350 5150
rect -250 5050 -200 5150
rect -550 4200 -200 5050
rect -550 4100 -350 4200
rect -250 4100 -200 4200
rect -550 3250 -200 4100
rect -550 3150 -350 3250
rect -250 3150 -200 3250
rect -550 2300 -200 3150
rect -550 2200 -350 2300
rect -250 2200 -200 2300
rect -550 1350 -200 2200
rect 3050 7050 3450 7200
rect 3050 6350 3100 7050
rect 3150 6350 3450 7050
rect 3050 6100 3450 6350
rect 3050 5400 3100 6100
rect 3150 5400 3450 6100
rect 3050 5150 3450 5400
rect 3050 4450 3100 5150
rect 3150 4450 3450 5150
rect 3050 4200 3450 4450
rect 3050 3500 3100 4200
rect 3150 3500 3450 4200
rect 3050 3250 3450 3500
rect 3050 2550 3100 3250
rect 3150 2550 3450 3250
rect 3050 2300 3450 2550
rect 3050 1600 3100 2300
rect 3150 1600 3450 2300
rect 3050 1500 3450 1600
rect -550 1250 -350 1350
rect -250 1250 -200 1350
rect -550 500 -200 1250
rect -650 -400 3550 500
<< labels >>
rlabel locali -650 650 -650 650 3 D6
port 2 e
rlabel locali -650 1600 -650 1600 3 D5
port 3 e
rlabel locali -650 2550 -650 2550 3 D4
port 4 e
rlabel locali -650 3500 -650 3500 3 D3
port 5 e
rlabel locali -650 4450 -650 4450 3 D2
port 6 e
rlabel locali -650 5400 -650 5400 3 D1
port 7 e
rlabel locali -650 6350 -650 6350 3 D0
port 8 e
rlabel locali -650 8600 -650 8600 3 Vc
port 9 e
rlabel locali -650 8800 -650 8800 3 Vg
port 10 e
rlabel metal1 -650 50 -650 50 3 GND
port 11 e
rlabel locali -650 8400 -650 8400 3 Vbn
port 12 e
rlabel metal1 -650 7650 -650 7650 3 VDD
port 13 e
rlabel locali 3550 -550 3550 -550 3 Iout
port 1 e
<< end >>
