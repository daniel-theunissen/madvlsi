magic
tech sky130A
timestamp 1762129613
<< nwell >>
rect -350 1800 950 3700
<< nmos >>
rect 0 1250 400 1550
rect 0 800 400 1100
rect 0 350 400 650
rect 0 -100 400 200
<< pmos >>
rect 0 3250 400 3550
rect 0 2800 400 3100
rect 0 2350 400 2650
rect 0 1900 400 2200
<< ndiff >>
rect -250 1450 0 1550
rect -250 1350 -150 1450
rect -100 1350 0 1450
rect -250 1250 0 1350
rect 400 1450 650 1550
rect 400 1350 500 1450
rect 550 1350 650 1450
rect 400 1250 650 1350
rect -250 1000 0 1100
rect -250 900 -150 1000
rect -100 900 0 1000
rect -250 800 0 900
rect 400 1000 650 1100
rect 400 900 500 1000
rect 550 900 650 1000
rect 400 800 650 900
rect -250 550 0 650
rect -250 450 -150 550
rect -100 450 0 550
rect -250 350 0 450
rect 400 550 650 650
rect 400 450 500 550
rect 550 450 650 550
rect 400 350 650 450
rect -250 100 0 200
rect -250 0 -150 100
rect -100 0 0 100
rect -250 -100 0 0
rect 400 100 650 200
rect 400 0 500 100
rect 550 0 650 100
rect 400 -100 650 0
<< pdiff >>
rect -250 3450 0 3550
rect -250 3350 -150 3450
rect -100 3350 0 3450
rect -250 3250 0 3350
rect 400 3450 650 3550
rect 400 3350 500 3450
rect 550 3350 650 3450
rect 400 3250 650 3350
rect -250 3000 0 3100
rect -250 2900 -150 3000
rect -100 2900 0 3000
rect -250 2800 0 2900
rect 400 3000 650 3100
rect 400 2900 500 3000
rect 550 2900 650 3000
rect 400 2800 650 2900
rect -250 2550 0 2650
rect -250 2450 -150 2550
rect -100 2450 0 2550
rect -250 2350 0 2450
rect 400 2550 650 2650
rect 400 2450 500 2550
rect 550 2450 650 2550
rect 400 2350 650 2450
rect -250 2100 0 2200
rect -250 2000 -150 2100
rect -100 2000 0 2100
rect -250 1900 0 2000
rect 400 2100 650 2200
rect 400 2000 500 2100
rect 550 2000 650 2100
rect 400 1900 650 2000
<< ndiffc >>
rect -150 1350 -100 1450
rect 500 1350 550 1450
rect -150 900 -100 1000
rect 500 900 550 1000
rect -150 450 -100 550
rect 500 450 550 550
rect -150 0 -100 100
rect 500 0 550 100
<< pdiffc >>
rect -150 3350 -100 3450
rect 500 3350 550 3450
rect -150 2900 -100 3000
rect 500 2900 550 3000
rect -150 2450 -100 2550
rect 500 2450 550 2550
rect -150 2000 -100 2100
rect 500 2000 550 2100
<< psubdiff >>
rect -500 550 -250 650
rect -500 450 -400 550
rect -350 450 -250 550
rect -500 350 -250 450
<< nsubdiff >>
rect 650 3000 900 3100
rect 650 2900 750 3000
rect 800 2900 900 3000
rect 650 2800 900 2900
<< psubdiffcont >>
rect -400 450 -350 550
<< nsubdiffcont >>
rect 750 2900 800 3000
<< poly >>
rect 0 3650 400 3700
rect 0 3600 50 3650
rect 350 3600 400 3650
rect 0 3550 400 3600
rect 0 3100 400 3250
rect 0 2650 400 2800
rect 0 2200 400 2350
rect 0 1850 400 1900
rect 0 1650 400 1700
rect 0 1600 50 1650
rect 350 1600 400 1650
rect 0 1550 400 1600
rect 0 1200 400 1250
rect 0 1100 400 1150
rect 0 650 400 800
rect 0 200 400 350
rect 0 -150 400 -100
rect 0 -200 50 -150
rect 350 -200 400 -150
rect 0 -250 400 -200
<< polycont >>
rect 50 3600 350 3650
rect 50 1600 350 1650
rect 50 -200 350 -150
<< locali >>
rect -550 3700 400 3750
rect -550 3600 -100 3650
rect 0 3600 50 3650
rect 350 3600 400 3700
rect -150 3500 -100 3600
rect -200 3450 -50 3500
rect -200 3350 -150 3450
rect -100 3350 -50 3450
rect -300 3300 -50 3350
rect 450 3450 600 3500
rect 450 3350 500 3450
rect 550 3350 600 3450
rect 450 3300 600 3350
rect -300 1650 -250 3300
rect 500 3050 550 3300
rect -200 3000 -50 3050
rect -200 2900 -150 3000
rect -100 2900 -50 3000
rect -200 2850 -50 2900
rect 450 3000 600 3050
rect 450 2900 500 3000
rect 550 2900 600 3000
rect 450 2850 600 2900
rect 700 3000 850 3050
rect 700 2900 750 3000
rect 800 2900 850 3000
rect 700 2850 850 2900
rect -150 2600 -100 2850
rect -200 2550 -50 2600
rect -200 2450 -150 2550
rect -100 2450 -50 2550
rect -200 2400 -50 2450
rect 450 2550 600 2600
rect 450 2450 500 2550
rect 550 2450 600 2550
rect 450 2400 600 2450
rect 500 2150 550 2400
rect -200 2100 -50 2150
rect -200 2000 -150 2100
rect -100 2000 -50 2100
rect -200 1950 -50 2000
rect 450 2100 600 2150
rect 450 2000 500 2100
rect 550 2000 600 2100
rect 450 1950 600 2000
rect -150 1800 -100 1950
rect -150 1750 700 1800
rect -300 1600 50 1650
rect 350 1600 400 1650
rect -150 1500 -100 1600
rect -200 1450 -50 1500
rect -200 1350 -150 1450
rect -100 1350 -50 1450
rect -200 1300 -50 1350
rect 450 1450 600 1500
rect 450 1350 500 1450
rect 550 1350 600 1450
rect 450 1300 600 1350
rect 500 1050 550 1300
rect -200 1000 -50 1050
rect -200 900 -150 1000
rect -100 900 -50 1000
rect -200 850 -50 900
rect 450 1000 600 1050
rect 450 900 500 1000
rect 550 900 600 1000
rect 450 850 600 900
rect 500 600 550 850
rect -450 550 -300 600
rect -450 450 -400 550
rect -350 450 -300 550
rect -450 400 -300 450
rect -200 550 -50 600
rect -200 450 -150 550
rect -100 450 -50 550
rect -200 400 -50 450
rect 450 550 600 600
rect 450 450 500 550
rect 550 450 600 550
rect 450 400 600 450
rect -150 150 -100 400
rect 500 150 550 400
rect -200 100 -50 150
rect -200 0 -150 100
rect -100 0 -50 100
rect -200 -50 -50 0
rect 450 100 600 150
rect 450 0 500 100
rect 550 0 600 100
rect 450 -50 600 0
rect -150 -150 -100 -50
rect 650 -150 700 1750
rect -150 -200 50 -150
rect 350 -200 700 -150
<< viali >>
rect 500 3350 550 3450
rect 750 2900 800 3000
rect -150 900 -100 1000
rect -400 450 -350 550
<< metal1 >>
rect -550 3450 1000 3550
rect -550 3350 500 3450
rect 550 3350 1000 3450
rect -550 3250 1000 3350
rect 700 3000 850 3250
rect 700 2900 750 3000
rect 800 2900 850 3000
rect 700 2850 850 2900
rect -200 1000 -50 1050
rect -200 900 -150 1000
rect -100 900 -50 1000
rect -450 550 -300 600
rect -450 450 -400 550
rect -350 450 -300 550
rect -450 200 -300 450
rect -200 200 -50 900
rect -550 -100 1000 200
<< labels >>
rlabel locali -550 3725 -550 3725 7 Vbp
port 1 w
rlabel metal1 -550 3400 -550 3400 7 VDD
port 2 w
rlabel locali -550 3625 -550 3625 7 Vc
port 3 w
rlabel metal1 -550 50 -550 50 7 GND
port 4 w
<< end >>
