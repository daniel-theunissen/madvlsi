magic
tech sky130A
timestamp 1762026219
<< error_p >>
rect -150 -300 -100 -250
rect 200 -300 250 -250
rect 550 -300 600 -250
rect 900 -300 950 -250
rect 1250 -300 1300 -250
rect 1600 -300 1650 -250
rect 1950 -300 2000 -250
rect -250 -450 50 -300
rect 100 -450 400 -300
rect 450 -450 750 -300
rect 800 -450 1100 -300
rect 1150 -450 1450 -300
rect 1500 -450 1800 -300
rect 1850 -450 2150 -300
rect -250 -1000 50 -850
rect 100 -1000 400 -850
rect 450 -1000 750 -850
rect 800 -1000 1100 -850
rect 1150 -1000 1450 -850
rect 1500 -1000 1800 -850
rect 1850 -1000 2150 -850
rect -250 -1550 50 -1400
rect 100 -1550 400 -1400
rect 450 -1550 750 -1400
rect 800 -1550 1100 -1400
rect 1150 -1550 1450 -1400
rect 1500 -1550 1800 -1400
rect 1850 -1550 2150 -1400
<< nmos >>
rect -300 2650 600 2850
rect 650 2650 1550 2850
rect 1600 2650 2500 2850
rect 2550 2650 3450 2850
rect 3500 2650 4400 2850
rect 4450 2650 5350 2850
rect 5400 2650 6300 2850
rect 6350 2650 7250 2850
rect 7300 2650 8200 2850
rect 650 2150 1550 2350
rect 1600 2150 2500 2350
rect 2550 2150 3450 2350
rect 3500 2150 4400 2350
rect 4450 2150 5350 2350
rect 5400 2150 6300 2350
rect 650 1700 1550 1900
rect 1600 1700 2500 1900
rect 2550 1700 3450 1900
rect 3500 1700 4400 1900
rect 4450 1700 5350 1900
rect 5400 1700 6300 1900
rect -150 -250 -100 150
rect 200 -250 250 150
rect 550 -250 600 150
rect 900 -250 950 150
rect 1250 -250 1300 150
rect 1600 -250 1650 150
rect 1950 -250 2000 150
rect -250 -850 50 -450
rect 100 -850 400 -450
rect 450 -850 750 -450
rect 800 -850 1100 -450
rect 1150 -850 1450 -450
rect 1500 -850 1800 -450
rect 1850 -850 2150 -450
rect -250 -1400 50 -1000
rect 100 -1400 400 -1000
rect 450 -1400 750 -1000
rect 800 -1400 1100 -1000
rect 1150 -1400 1450 -1000
rect 1500 -1400 1800 -1000
rect 1850 -1400 2150 -1000
<< ndiff >>
rect -300 3000 600 3100
rect -300 2950 -200 3000
rect 500 2950 600 3000
rect -300 2850 600 2950
rect 650 3000 1550 3100
rect 650 2950 750 3000
rect 1450 2950 1550 3000
rect 650 2850 1550 2950
rect 1600 3000 2500 3100
rect 1600 2950 1700 3000
rect 2400 2950 2500 3000
rect 1600 2850 2500 2950
rect 2550 3000 3450 3100
rect 2550 2950 2650 3000
rect 3350 2950 3450 3000
rect 2550 2850 3450 2950
rect 3500 3000 4400 3100
rect 3500 2950 3600 3000
rect 4300 2950 4400 3000
rect 3500 2850 4400 2950
rect 4450 3000 5350 3100
rect 4450 2950 4550 3000
rect 5250 2950 5350 3000
rect 4450 2850 5350 2950
rect 5400 3000 6300 3100
rect 5400 2950 5500 3000
rect 6200 2950 6300 3000
rect 5400 2850 6300 2950
rect 6350 3000 7250 3100
rect 6350 2950 6450 3000
rect 7150 2950 7250 3000
rect 6350 2850 7250 2950
rect 7300 3000 8200 3100
rect 7300 2950 7400 3000
rect 8100 2950 8200 3000
rect 7300 2850 8200 2950
rect -300 2550 600 2650
rect -300 2500 -200 2550
rect 500 2500 600 2550
rect -300 2400 600 2500
rect 650 2550 1550 2650
rect 650 2500 750 2550
rect 1450 2500 1550 2550
rect 650 2350 1550 2500
rect 1600 2550 2500 2650
rect 1600 2500 1700 2550
rect 2400 2500 2500 2550
rect 1600 2350 2500 2500
rect 2550 2550 3450 2650
rect 2550 2500 2650 2550
rect 3350 2500 3450 2550
rect 2550 2350 3450 2500
rect 3500 2550 4400 2650
rect 3500 2500 3600 2550
rect 4300 2500 4400 2550
rect 3500 2350 4400 2500
rect 4450 2550 5350 2650
rect 4450 2500 4550 2550
rect 5250 2500 5350 2550
rect 4450 2350 5350 2500
rect 5400 2550 6300 2650
rect 5400 2500 5500 2550
rect 6200 2500 6300 2550
rect 5400 2350 6300 2500
rect 6350 2550 7250 2650
rect 6350 2500 6450 2550
rect 7150 2500 7250 2550
rect 6350 2400 7250 2500
rect 7300 2550 8200 2650
rect 7300 2500 7400 2550
rect 8100 2500 8200 2550
rect 7300 2400 8200 2500
rect 650 2050 1550 2150
rect 650 2000 750 2050
rect 1450 2000 1550 2050
rect 650 1900 1550 2000
rect 1600 2050 2500 2150
rect 1600 2000 1700 2050
rect 2400 2000 2500 2050
rect 1600 1900 2500 2000
rect 2550 2050 3450 2150
rect 2550 2000 3050 2050
rect 3350 2000 3450 2050
rect 2550 1900 3450 2000
rect 3500 2050 4400 2150
rect 3500 2000 4050 2050
rect 4350 2000 4400 2050
rect 3500 1900 4400 2000
rect 4450 2050 5350 2150
rect 4450 2000 4550 2050
rect 5250 2000 5350 2050
rect 4450 1900 5350 2000
rect 5400 2050 6300 2150
rect 5400 2000 5500 2050
rect 6200 2000 6300 2050
rect 5400 1900 6300 2000
rect 650 1600 1550 1700
rect 650 1550 750 1600
rect 1450 1550 1550 1600
rect 650 1450 1550 1550
rect 1600 1600 2500 1700
rect 1600 1550 1700 1600
rect 2400 1550 2500 1600
rect 1600 1450 2500 1550
rect 2550 1600 3450 1700
rect 2550 1550 2650 1600
rect 3350 1550 3450 1600
rect 2550 1450 3450 1550
rect 3500 1600 4400 1700
rect 3500 1550 3600 1600
rect 4300 1550 4400 1600
rect 3500 1450 4400 1550
rect 4450 1600 5350 1700
rect 4450 1550 4550 1600
rect 5250 1550 5350 1600
rect 4450 1450 5350 1550
rect 5400 1600 6300 1700
rect 5400 1550 5500 1600
rect 6200 1550 6300 1600
rect 5400 1450 6300 1550
rect -150 150 -100 200
rect 200 150 250 200
rect 550 150 600 200
rect 900 150 950 200
rect 1250 150 1300 200
rect 1600 150 1650 200
rect 1950 150 2000 200
rect -150 -300 -100 -250
rect 200 -300 250 -250
rect 550 -300 600 -250
rect 900 -300 950 -250
rect 1250 -300 1300 -250
rect 1600 -300 1650 -250
rect 1950 -300 2000 -250
rect -250 -450 50 -300
rect 100 -450 400 -300
rect 450 -450 750 -300
rect 800 -450 1100 -300
rect 1150 -450 1450 -300
rect 1500 -450 1800 -300
rect 1850 -450 2150 -300
rect -250 -1000 50 -850
rect 100 -1000 400 -850
rect 450 -1000 750 -850
rect 800 -1000 1100 -850
rect 1150 -1000 1450 -850
rect 1500 -1000 1800 -850
rect 1850 -1000 2150 -850
rect -250 -1550 50 -1400
rect 100 -1550 400 -1400
rect 450 -1550 750 -1400
rect 800 -1550 1100 -1400
rect 1150 -1550 1450 -1400
rect 1500 -1550 1800 -1400
rect 1850 -1550 2150 -1400
<< ndiffc >>
rect -200 2950 500 3000
rect 750 2950 1450 3000
rect 1700 2950 2400 3000
rect 2650 2950 3350 3000
rect 3600 2950 4300 3000
rect 4550 2950 5250 3000
rect 5500 2950 6200 3000
rect 6450 2950 7150 3000
rect 7400 2950 8100 3000
rect -200 2500 500 2550
rect 750 2500 1450 2550
rect 1700 2500 2400 2550
rect 2650 2500 3350 2550
rect 3600 2500 4300 2550
rect 4550 2500 5250 2550
rect 5500 2500 6200 2550
rect 6450 2500 7150 2550
rect 7400 2500 8100 2550
rect 750 2000 1450 2050
rect 1700 2000 2400 2050
rect 3050 2000 3350 2050
rect 4050 2000 4350 2050
rect 4550 2000 5250 2050
rect 5500 2000 6200 2050
rect 750 1550 1450 1600
rect 1700 1550 2400 1600
rect 2650 1550 3350 1600
rect 3600 1550 4300 1600
rect 4550 1550 5250 1600
rect 5500 1550 6200 1600
<< psubdiff >>
rect -300 3250 600 3350
rect -300 3200 -200 3250
rect 500 3200 600 3250
rect -300 3100 600 3200
rect 1600 3250 2500 3350
rect 1600 3200 1700 3250
rect 2400 3200 2500 3250
rect 1600 3100 2500 3200
rect 3500 3250 4400 3350
rect 3500 3200 3600 3250
rect 4300 3200 4400 3250
rect 3500 3100 4400 3200
rect 5400 3250 6300 3350
rect 5400 3200 5500 3250
rect 6200 3200 6300 3250
rect 5400 3100 6300 3200
rect 7300 3250 8200 3350
rect 7300 3200 7400 3250
rect 8100 3200 8200 3250
rect 7300 3100 8200 3200
rect 650 1350 1550 1450
rect 650 1300 750 1350
rect 1450 1300 1550 1350
rect 650 1200 1550 1300
rect 1600 1350 2500 1450
rect 1600 1300 1700 1350
rect 2400 1300 2500 1350
rect 1600 1200 2500 1300
rect 2550 1350 3450 1450
rect 2550 1300 2650 1350
rect 3350 1300 3450 1350
rect 2550 1200 3450 1300
rect 3500 1350 4400 1450
rect 3500 1300 3600 1350
rect 4300 1300 4400 1350
rect 3500 1200 4400 1300
rect 4450 1350 5350 1450
rect 4450 1300 4550 1350
rect 5250 1300 5350 1350
rect 4450 1200 5350 1300
rect 5400 1350 6300 1450
rect 5400 1300 5500 1350
rect 6200 1300 6300 1350
rect 5400 1200 6300 1300
<< psubdiffcont >>
rect -200 3200 500 3250
rect 1700 3200 2400 3250
rect 3600 3200 4300 3250
rect 5500 3200 6200 3250
rect 7400 3200 8100 3250
rect 750 1300 1450 1350
rect 1700 1300 2400 1350
rect 2650 1300 3350 1350
rect 3600 1300 4300 1350
rect 4550 1300 5250 1350
rect 5500 1300 6200 1350
<< poly >>
rect -450 2650 -300 2850
rect 600 2650 650 2850
rect 1550 2650 1600 2850
rect 2500 2650 2550 2850
rect 3450 2650 3500 2850
rect 4400 2650 4450 2850
rect 5350 2650 5400 2850
rect 6300 2650 6350 2850
rect 7250 2650 7300 2850
rect 8200 2650 8350 2850
rect -450 2150 650 2350
rect 1550 2150 1600 2350
rect 2500 2150 2550 2350
rect 3450 2150 3500 2350
rect 4400 2150 4450 2350
rect 5350 2150 5400 2350
rect 6300 2150 8350 2350
rect -450 1700 650 1900
rect 1550 1700 1600 1900
rect 2500 1700 2550 1900
rect 3450 1700 3500 1900
rect 4400 1700 4450 1900
rect 5350 1700 5400 1900
rect 6300 1700 8350 1900
rect -250 -250 -150 150
rect -100 -250 50 150
rect 100 -250 200 150
rect 250 -250 400 150
rect 450 -250 550 150
rect 600 -250 750 150
rect 800 -250 900 150
rect 950 -250 1100 150
rect 1150 -250 1250 150
rect 1300 -250 1450 150
rect 1500 -250 1600 150
rect 1650 -250 1800 150
rect 1850 -250 1950 150
rect 2000 -250 2150 150
rect -400 -850 -250 -450
rect 50 -850 100 -450
rect 400 -850 450 -450
rect 750 -850 800 -450
rect 1100 -850 1150 -450
rect 1450 -850 1500 -450
rect 1800 -850 1850 -450
rect 2150 -850 2300 -450
rect -400 -1400 -250 -1000
rect 50 -1400 100 -1000
rect 400 -1400 450 -1000
rect 750 -1400 800 -1000
rect 1100 -1400 1150 -1000
rect 1450 -1400 1500 -1000
rect 1800 -1400 1850 -1000
rect 2150 -1400 2300 -1000
<< locali >>
rect -250 3250 550 3300
rect -250 3200 -200 3250
rect 500 3200 550 3250
rect -250 3050 550 3200
rect 1650 3250 2450 3300
rect 1650 3200 1700 3250
rect 2400 3200 2450 3250
rect 1650 3050 2450 3200
rect 3550 3250 4350 3300
rect 3550 3200 3600 3250
rect 4300 3200 4350 3250
rect 3550 3050 4350 3200
rect 5450 3250 6250 3300
rect 5450 3200 5500 3250
rect 6200 3200 6250 3250
rect 5450 3050 6250 3200
rect 7350 3250 8150 3300
rect 7350 3200 7400 3250
rect 8100 3200 8150 3250
rect 7350 3050 8150 3200
rect -250 3000 6250 3050
rect -250 2950 -200 3000
rect 500 2950 750 3000
rect 1450 2950 1700 3000
rect 2400 2950 2650 3000
rect 3350 2950 3600 3000
rect 4300 2950 4550 3000
rect 5250 2950 5500 3000
rect 6200 2950 6250 3000
rect -250 2900 6250 2950
rect 6400 3000 8150 3050
rect 6400 2950 6450 3000
rect 7150 2950 7400 3000
rect 8100 2950 8150 3000
rect 6400 2900 8150 2950
rect -250 2550 1500 2600
rect -250 2500 -200 2550
rect 500 2500 750 2550
rect 1450 2500 1500 2550
rect -250 2450 1500 2500
rect 1650 2550 2450 2600
rect 1650 2500 1700 2550
rect 2400 2500 2450 2550
rect 1650 2450 2450 2500
rect 2600 2550 3400 2600
rect 2600 2500 2650 2550
rect 3350 2500 3400 2550
rect 2600 2450 3400 2500
rect 3550 2550 4350 2600
rect 3550 2500 3600 2550
rect 4300 2500 4350 2550
rect 3550 2450 4350 2500
rect 4500 2550 5300 2600
rect 4500 2500 4550 2550
rect 5250 2500 5300 2550
rect 4500 2450 5300 2500
rect 5450 2550 6250 2600
rect 5450 2500 5500 2550
rect 6200 2500 6250 2550
rect 5450 2450 6250 2500
rect 6400 2550 8150 2600
rect 6400 2500 6450 2550
rect 7150 2500 7400 2550
rect 8100 2500 8150 2550
rect 6400 2450 8150 2500
rect 700 2050 1550 2100
rect 700 2000 750 2050
rect 1450 2000 1550 2050
rect 700 1950 1550 2000
rect 1650 2050 2500 2100
rect 1650 2000 1700 2050
rect 2400 2000 2500 2050
rect 1650 1950 2500 2000
rect 3050 2050 3450 2100
rect 3350 2000 3450 2050
rect 3050 1950 3450 2000
rect 4000 2050 4350 2100
rect 4000 2000 4050 2050
rect 4000 1950 4350 2000
rect 4500 2050 5350 2100
rect 4500 2000 4550 2050
rect 5250 2000 5350 2050
rect 4500 1950 5350 2000
rect 5450 2050 6300 2100
rect 5450 2000 5500 2050
rect 6200 2000 6300 2050
rect 5450 1950 6300 2000
rect 700 1600 1500 1650
rect 700 1550 750 1600
rect 1450 1550 1500 1600
rect 700 1350 1500 1550
rect 700 1300 750 1350
rect 1450 1300 1500 1350
rect 700 1250 1500 1300
rect 1650 1600 2450 1650
rect 1650 1550 1700 1600
rect 2400 1550 2450 1600
rect 1650 1350 2450 1550
rect 1650 1300 1700 1350
rect 2400 1300 2450 1350
rect 1650 1250 2450 1300
rect 2600 1600 3400 1650
rect 2600 1550 2650 1600
rect 3350 1550 3400 1600
rect 2600 1350 3400 1550
rect 2600 1300 2650 1350
rect 3350 1300 3400 1350
rect 2600 1250 3400 1300
rect 3550 1600 4350 1650
rect 3550 1550 3600 1600
rect 4300 1550 4350 1600
rect 3550 1350 4350 1550
rect 3550 1300 3600 1350
rect 4300 1300 4350 1350
rect 3550 1250 4350 1300
rect 4500 1600 5300 1650
rect 4500 1550 4550 1600
rect 5250 1550 5300 1600
rect 4500 1350 5300 1550
rect 4500 1300 4550 1350
rect 5250 1300 5300 1350
rect 4500 1250 5300 1300
rect 5450 1600 6250 1650
rect 5450 1550 5500 1600
rect 6200 1550 6250 1600
rect 5450 1350 6250 1550
rect 5450 1300 5500 1350
rect 6200 1300 6250 1350
rect 5450 1250 6250 1300
<< end >>
