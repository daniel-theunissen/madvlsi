* SPICE3 file created from mirror.ext - technology: sky130A

.subckt mirror Iin Iout Vbn VDD GND
X0 a_1220_n60# Vbn a_570_n60# GND sky130_fd_pr__nfet_01v8 ad=0.375 pd=3.25 as=0.375 ps=3.25 w=3 l=3
X1 a_n30_660# Vbn a_1220_n60# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.375 ps=3.25 w=3 l=3
X2 VDD a_n940_n770# a_n180_1480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=3
X3 a_n30_660# a_n30_660# a_n130_690# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=3
X4 a_3740_1450# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X5 a_2880_1450# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X6 a_n130_690# a_n950_440# a_n950_440# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X7 GND Vbn a_5040_n60# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0.375 ps=3.25 w=3 l=3
X8 Iin a_3740_1450# a_2880_1450# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X9 a_3570_440# a_3570_440# a_4290_690# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=3
X10 a_n940_n770# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X11 a_570_n60# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=0.375 pd=3.25 as=0.75 ps=3.5 w=3 l=3
X12 GND Vbn a_n950_440# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X13 a_3480_1480# a_4440_1450# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=3
X14 a_5040_n60# Vbn a_4390_n60# GND sky130_fd_pr__nfet_01v8 ad=0.375 pd=3.25 as=0.375 ps=3.25 w=3 l=3
X15 a_n130_690# a_n30_660# a_n30_660# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=3
X16 VDD a_n30_660# a_n130_690# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X17 GND Vbn a_620_n770# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X18 GND Vbn a_2880_1450# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X19 GND Vbn a_4440_1450# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X20 a_n180_1480# a_n950_440# a_n940_n770# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X21 Iout a_620_n770# a_n180_1480# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X22 a_4390_n60# Vbn a_3570_440# GND sky130_fd_pr__nfet_01v8 ad=0.375 pd=3.25 as=1.5 ps=7 w=3 l=3
X23 GND Vbn a_n940_n770# GND sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X24 a_4290_690# a_3570_440# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=1.5 ps=7 w=3 l=3
X25 Iin a_n940_n770# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=3
X26 a_4440_1450# a_3740_1450# a_3480_1480# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X27 a_620_n770# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X28 a_4440_1450# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X29 VDD a_4440_1450# Iin VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=3
X30 a_3740_1450# a_3740_1450# a_4290_690# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X31 a_3480_1480# a_2880_1450# Iout VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
X32 a_4290_690# a_3570_440# a_3570_440# VDD sky130_fd_pr__pfet_01v8 ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=3
X33 a_620_n770# a_n950_440# Iin VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=7 as=0.75 ps=3.5 w=3 l=3
.ends

