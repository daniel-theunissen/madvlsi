* SPICE3 file created from mag_cascode_bias.ext - technology: sky130A

.subckt mag_cascode_bias Vbp VDD Vc GND
X0 a_800_n200# Vc Vc GND sky130_fd_pr__nfet_01v8 ad=7.5 pd=11 as=7.5 ps=11 w=3 l=4
X1 a_800_3800# Vbp a_n500_4700# VDD sky130_fd_pr__pfet_01v8 ad=7.5 pd=11 as=7.5 ps=11 w=3 l=4
X2 a_800_n200# a_n500_n200# a_n500_n200# GND sky130_fd_pr__nfet_01v8 ad=7.5 pd=11 as=7.5 ps=11 w=3 l=4
X3 VDD Vbp a_n500_4700# VDD sky130_fd_pr__pfet_01v8 ad=7.5 pd=11 as=7.5 ps=11 w=3 l=4
X4 VDD Vbp Vc VDD sky130_fd_pr__pfet_01v8 ad=7.5 pd=11 as=7.5 ps=11 w=3 l=4
X5 a_800_n200# a_n500_n200# a_n500_n200# GND sky130_fd_pr__nfet_01v8 ad=7.5 pd=11 as=7.5 ps=11 w=3 l=4
X6 a_800_n200# a_n500_n200# GND GND sky130_fd_pr__nfet_01v8 ad=7.5 pd=11 as=7.5 ps=11 w=3 l=4
X7 a_800_3800# Vbp a_n500_n200# VDD sky130_fd_pr__pfet_01v8 ad=7.5 pd=11 as=7.5 ps=11 w=3 l=4
.ends

