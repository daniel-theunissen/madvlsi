magic
tech sky130A
timestamp 1762122893
<< error_p >>
rect -750 5200 -450 5500
rect -50 5200 250 5500
rect -750 4600 -450 4900
rect -50 4600 250 4900
rect -1500 4000 -1200 4300
rect -800 4000 -450 4300
rect -50 4000 250 4300
rect -750 3400 -450 3700
rect -50 3400 250 3700
rect -1500 2800 -1200 3100
rect -800 2800 -450 3100
rect -50 2800 250 3100
rect -750 2200 -450 2500
rect -50 2200 250 2500
rect -1500 1600 -1200 1900
rect -800 1600 -450 1900
rect -50 1600 250 1900
rect -1500 1000 -1200 1300
rect -800 1000 -450 1300
rect -50 1000 250 1300
<< nmos >>
rect -450 5200 -50 5500
rect -450 4600 -50 4900
rect -1200 4000 -800 4300
rect -450 4000 -50 4300
rect -450 3400 -50 3700
rect -1200 2800 -800 3100
rect -450 2800 -50 3100
rect -450 2200 -50 2500
rect -1200 1600 -800 1900
rect -450 1600 -50 1900
rect -1200 1000 -800 1300
rect -450 1000 -50 1300
<< ndiff >>
rect -750 5200 -450 5500
rect -50 5200 250 5500
rect -750 4600 -450 4900
rect -50 4600 250 4900
rect -1500 4000 -1200 4300
rect -800 4000 -450 4300
rect -50 4000 250 4300
rect -750 3400 -450 3700
rect -50 3400 250 3700
rect -1500 2800 -1200 3100
rect -800 2800 -450 3100
rect -50 2800 250 3100
rect -750 2200 -450 2500
rect -50 2200 250 2500
rect -1500 1600 -1200 1900
rect -800 1600 -450 1900
rect -50 1600 250 1900
rect -1500 1000 -1200 1300
rect -800 1000 -450 1300
rect -50 1000 250 1300
<< poly >>
rect -1200 4300 -800 5650
rect -450 5500 -50 5650
rect -450 4900 -50 5200
rect -450 4300 -50 4600
rect -1200 3100 -800 4000
rect -450 3700 -50 4000
rect -450 3100 -50 3400
rect -1200 1900 -800 2800
rect -450 2500 -50 2800
rect -450 1900 -50 2200
rect -1200 1300 -800 1600
rect -450 1300 -50 1600
rect -1200 850 -800 1000
rect -450 850 -50 1000
<< end >>
