* SPICE3 file created from mag_current_div.ext - technology: sky130A

.subckt mag_current_div Vbp VDD Vbn2 GND
X0 a_n6100_9200# Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=6 ps=10 w=3 l=4
X1 a_n2400_8000# GND a_n2400_5600# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=3.75 ps=5.5 w=3 l=4
X2 Vbn2 Vbn2 GND GND sky130_fd_pr__nfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=3
X3 a_n2400_11600# GND a_n2400_10400# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=6 ps=10 w=3 l=4
X4 a_n4900_2000# GND a_n6100_2000# VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=6 ps=10 w=3 l=4
X5 a_n6100_2000# GND a_n6100_4400# VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=6 ps=10 w=3 l=4
X6 a_n2400_11600# GND GND VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=3 ps=5 w=3 l=4
X7 a_n2400_11600# GND a_n2400_10400# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=3.75 ps=5.5 w=3 l=4
X8 a_n6100_6800# GND a_n6100_9200# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=6 ps=10 w=3 l=4
X9 Vbn2 GND a_n4900_2000# VDD sky130_fd_pr__pfet_01v8 ad=3 pd=5 as=3.75 ps=5.5 w=3 l=4
X10 GND Vbn2 Vbn2 GND sky130_fd_pr__nfet_01v8 ad=6 pd=10 as=3 ps=5 w=3 l=3
X11 GND GND a_n6100_9200# VDD sky130_fd_pr__pfet_01v8 ad=3 pd=5 as=3.75 ps=5.5 w=3 l=4
X12 a_n6100_6800# GND a_n6100_9200# VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=6 ps=10 w=3 l=4
X13 a_n2400_8000# GND GND VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=3 ps=5 w=3 l=4
X14 a_n2400_5600# GND a_n2400_2000# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=3.75 ps=5.5 w=3 l=4
X15 a_n2400_10400# GND a_n2400_8000# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=6 ps=10 w=3 l=4
X16 a_n4900_2000# GND a_n6100_2000# VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=6 ps=10 w=3 l=4
X17 a_n6100_4400# GND a_n6100_6800# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=6 ps=10 w=3 l=4
X18 a_n2400_2000# GND Vbn2 VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=3 ps=5 w=3 l=4
X19 a_n2400_11600# GND GND VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=3 ps=5 w=3 l=4
X20 a_n2400_5600# GND GND VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=3 ps=5 w=3 l=4
X21 GND GND a_n6100_6800# VDD sky130_fd_pr__pfet_01v8 ad=3 pd=5 as=3.75 ps=5.5 w=3 l=4
X22 a_n2400_8000# GND a_n2400_5600# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=6 ps=10 w=3 l=4
X23 GND GND a_n6100_4400# VDD sky130_fd_pr__pfet_01v8 ad=3 pd=5 as=3.75 ps=5.5 w=3 l=4
X24 a_n2400_10400# GND a_n2400_8000# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=3.75 ps=5.5 w=3 l=4
X25 a_n2400_10400# GND GND VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=3 ps=5 w=3 l=4
X26 a_n6100_2000# GND a_n6100_4400# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=6 ps=10 w=3 l=4
X27 a_n2400_2000# GND Vbn2 VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=3 ps=5 w=3 l=4
X28 a_n6100_4400# GND a_n6100_6800# VDD sky130_fd_pr__pfet_01v8 ad=3.75 pd=5.5 as=6 ps=10 w=3 l=4
X29 VDD Vbp a_n2400_11600# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=3.75 ps=5.5 w=3 l=4
X30 Vbn2 GND a_n4900_2000# VDD sky130_fd_pr__pfet_01v8 ad=3 pd=5 as=3.75 ps=5.5 w=3 l=4
X31 GND GND a_n6100_9200# VDD sky130_fd_pr__pfet_01v8 ad=3 pd=5 as=6 ps=10 w=3 l=4
X32 GND GND a_n6100_2000# VDD sky130_fd_pr__pfet_01v8 ad=3 pd=5 as=3.75 ps=5.5 w=3 l=4
X33 a_n2400_5600# GND a_n2400_2000# VDD sky130_fd_pr__pfet_01v8 ad=6 pd=10 as=3.75 ps=5.5 w=3 l=4
.ends

