* NGSPICE file created from controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

.subckt controller GND VDD ADC0 ADC1 ADC2 ADC3 ADC4
+ ADC5 ADC6 ADC7 clk comp DAC0 DAC1 DAC2 DAC3
+ DAC4 DAC5 DAC6 DAC7 rst_n
XFILLER_3_89 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_66 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_062_ net2 _029_ GND GND VDD VDD _030_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_165 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_114_ clknet_1_1__leaf_clk _010_ GND GND VDD VDD net3 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_35 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput7 net7 GND GND VDD VDD ADC4 sky130_fd_sc_hd__buf_2
XFILLER_9_138 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_3_57 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_67 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_14 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_69 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_061_ net20 count\[0\] count\[2\] net19 GND GND VDD VDD _029_ sky130_fd_sc_hd__or4b_2
X_113_ clknet_1_1__leaf_clk _009_ GND GND VDD VDD net16 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_225 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_253 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_36 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput8 net8 GND GND VDD VDD ADC5 sky130_fd_sc_hd__buf_2
Xoutput10 net10 GND GND VDD VDD ADC7 sky130_fd_sc_hd__buf_2
XFILLER_3_69 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_68 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_131 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_13 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_060_ net20 net21 count\[2\] GND GND VDD VDD _028_ sky130_fd_sc_hd__nor3_1
XFILLER_9_57 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_112_ clknet_1_0__leaf_clk _008_ GND GND VDD VDD net15 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_215 GND GND VDD VDD sky130_fd_sc_hd__decap_8
Xhold10 _016_ GND GND VDD VDD net31 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput11 net11 GND GND VDD VDD DAC0 sky130_fd_sc_hd__buf_2
XFILLER_0_221 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_37 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput9 net9 GND GND VDD VDD ADC6 sky130_fd_sc_hd__buf_2
XFILLER_8_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_3_15 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_7 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_69 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_121 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_5_143 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_9_69 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_47 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_9_25 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_111_ clknet_1_0__leaf_clk _007_ GND GND VDD VDD net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_81 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xhold11 net3 GND GND VDD VDD net32 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_15 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xoutput12 net12 GND GND VDD VDD DAC1 sky130_fd_sc_hd__buf_2
XFILLER_0_277 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_38 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_27 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_5_199 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_114 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_18 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xclkload0 clknet_1_0__leaf_clk GND GND VDD VDD clkload0/X sky130_fd_sc_hd__clkbuf_8
X_110_ clknet_1_0__leaf_clk _006_ GND GND VDD VDD net13 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_93 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xhold12 net6 GND GND VDD VDD net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
Xoutput13 net13 GND GND VDD VDD DAC2 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_39 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_39 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_197 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_153 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_5_167 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_29 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_126 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_9_281 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_70 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xhold13 _013_ GND GND VDD VDD net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_276 GND GND VDD VDD sky130_fd_sc_hd__decap_4
Xoutput14 net14 GND GND VDD VDD DAC3 sky130_fd_sc_hd__buf_2
XFILLER_5_113 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_71 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_099_ net18 net24 _049_ GND GND VDD VDD _017_ sky130_fd_sc_hd__mux2_1
XFILLER_1_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_29 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xoutput15 net15 GND GND VDD VDD DAC4 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_247 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_225 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_40 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_166 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_169 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_29 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_72 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_231 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_098_ net17 net30 _049_ GND GND VDD VDD _016_ sky130_fd_sc_hd__mux2_1
XFILLER_3_201 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_212 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xoutput16 net16 GND GND VDD VDD DAC5 sky130_fd_sc_hd__buf_2
XFILLER_0_237 GND GND VDD VDD sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk GND GND VDD VDD clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_7_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_8_189 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_41 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_41 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_170 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_73 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_20 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_243 GND GND VDD VDD sky130_fd_sc_hd__fill_1
X_097_ net16 net22 _049_ GND GND VDD VDD _015_ sky130_fd_sc_hd__mux2_1
Xoutput17 net17 GND GND VDD VDD DAC6 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_3_42 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_105 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_182 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_21 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_74 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_13 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_096_ net15 net27 _049_ GND GND VDD VDD _014_ sky130_fd_sc_hd__mux2_1
XFILLER_6_200 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_225 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xoutput18 net18 GND GND VDD VDD DAC7 sky130_fd_sc_hd__buf_2
X_079_ net20 net21 net19 count\[2\] GND GND VDD VDD _041_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_5_Right_5 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_43 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_158 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_7_180 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_4_65 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_194 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_1_142 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_22 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout20 count\[1\] GND GND VDD VDD net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_286 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_9_253 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_9_220 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_75 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_186 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_153 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
X_095_ net14 net33 _049_ GND GND VDD VDD _013_ sky130_fd_sc_hd__mux2_1
XFILLER_3_237 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_281 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_078_ _039_ _040_ _030_ GND GND VDD VDD _005_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_3_44 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xfanout21 count\[0\] GND GND VDD VDD net21 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_76 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_198 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_165 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_23 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_094_ net13 net26 _049_ GND GND VDD VDD _012_ sky130_fd_sc_hd__mux2_1
XFILLER_3_249 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_077_ net1 _023_ _037_ GND GND VDD VDD _040_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_55 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_7_77 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_141 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_233 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_77 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_24 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_093_ net12 net29 _049_ GND GND VDD VDD _011_ sky130_fd_sc_hd__mux2_1
XFILLER_6_269 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_1_57 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xinput1 comp GND GND VDD VDD net1 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_7_Left_17 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_076_ net20 net19 count\[2\] net21 GND GND VDD VDD _039_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_6_56 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_059_ net16 GND GND VDD VDD _027_ sky130_fd_sc_hd__inv_2
XFILLER_8_106 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_131 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_78 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_25 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_278 GND GND VDD VDD sky130_fd_sc_hd__fill_2
X_092_ net11 net32 _049_ GND GND VDD VDD _010_ sky130_fd_sc_hd__mux2_1
XFILLER_1_69 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xinput2 rst_n GND GND VDD VDD net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_281 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
X_075_ _036_ _038_ _030_ GND GND VDD VDD _004_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_6_57 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_57 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_058_ net15 GND GND VDD VDD _026_ sky130_fd_sc_hd__inv_2
XFILLER_8_118 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_7_140 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_121 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_26 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_146 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_1_113 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_79 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_15 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_091_ _021_ _029_ GND GND VDD VDD _049_ sky130_fd_sc_hd__or2_4
X_074_ net19 net1 _032_ _037_ GND GND VDD VDD _038_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_6_58 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_69 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_057_ net14 GND GND VDD VDD _025_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Right_0 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_109_ clknet_1_0__leaf_clk _005_ GND GND VDD VDD net12 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_185 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_15 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_27 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_125 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_9_225 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_9_203 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_1_169 GND GND VDD VDD sky130_fd_sc_hd__fill_1
X_090_ _047_ _048_ _030_ GND GND VDD VDD _009_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_27 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_59 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_073_ net21 net19 count\[2\] net20 GND GND VDD VDD _037_ sky130_fd_sc_hd__or4bb_1
XFILLER_7_15 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_056_ net13 GND GND VDD VDD _024_ sky130_fd_sc_hd__inv_2
X_108_ clknet_1_0__leaf_clk _004_ GND GND VDD VDD net11 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_197 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_9_248 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_28 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_81 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_39 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_262 GND GND VDD VDD sky130_fd_sc_hd__fill_1
X_072_ net19 _032_ net11 GND GND VDD VDD _036_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_221 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_055_ net12 GND GND VDD VDD _023_ sky130_fd_sc_hd__inv_2
XFILLER_7_27 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_107_ clknet_1_0__leaf_clk _003_ GND GND VDD VDD count\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_121 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_29 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_6_219 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_252 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_12 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_233 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_071_ _034_ _035_ _030_ GND GND VDD VDD _003_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_7_39 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_60 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_054_ net1 GND GND VDD VDD _022_ sky130_fd_sc_hd__inv_2
X_123_ clknet_1_1__leaf_clk _019_ GND GND VDD VDD net18 sky130_fd_sc_hd__dfxtp_1
X_106_ clknet_1_0__leaf_clk _002_ GND GND VDD VDD count\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_7_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_29 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_4_158 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_261 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_2_245 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_070_ net19 _032_ GND GND VDD VDD _035_ sky130_fd_sc_hd__nand2_1
XFILLER_4_3 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_122_ clknet_1_1__leaf_clk _018_ GND GND VDD VDD net17 sky130_fd_sc_hd__dfxtp_1
X_053_ net2 GND GND VDD VDD _021_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_61 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_105_ clknet_1_0__leaf_clk _001_ GND GND VDD VDD count\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_30 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_41 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_121_ clknet_1_1__leaf_clk net25 GND GND VDD VDD net10 sky130_fd_sc_hd__dfxtp_1
X_052_ net19 GND GND VDD VDD _020_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f_clk clknet_0_clk GND GND VDD VDD clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_7_62 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_104_ clknet_1_0__leaf_clk _000_ GND GND VDD VDD count\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 GND GND VDD VDD sky130_fd_sc_hd__decap_8
Xfanout19 count\[3\] GND GND VDD VDD net19 sky130_fd_sc_hd__buf_2
XFILLER_9_208 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_230 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_31 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_233 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_2_53 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_120_ clknet_1_1__leaf_clk net31 GND GND VDD VDD net9 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_6_Left_16 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_63 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_103_ _020_ _022_ _028_ _051_ _021_ GND GND VDD VDD _019_ sky130_fd_sc_hd__a311o_1
XFILLER_7_103 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_7_169 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_8_41 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_85 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_4_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xhold1 net8 GND GND VDD VDD net22 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_197 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_31 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_32 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_1_281 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_65 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_3 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_64 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_102_ _028_ net18 GND GND VDD VDD _051_ sky130_fd_sc_hd__and2b_1
XFILLER_6_181 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_8_53 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_151 GND GND VDD VDD sky130_fd_sc_hd__decap_8
Xhold2 _015_ GND GND VDD VDD net23 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_8_287 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_165 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_5_43 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_33 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_2_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_101_ _028_ _050_ net2 GND GND VDD VDD _018_ sky130_fd_sc_hd__o21a_1
XFILLER_6_193 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_8_65 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xhold3 net10 GND GND VDD VDD net24 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_34 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_225 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_100_ _022_ net17 _047_ GND GND VDD VDD _050_ sky130_fd_sc_hd__mux2_1
XFILLER_6_172 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_8_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_109 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xhold4 _017_ GND GND VDD VDD net25 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_45 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_201 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_0_3 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_162 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_8_89 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_46 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 net5 GND GND VDD VDD net26 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_11 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_9_193 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_6_141 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_089_ net1 _027_ _045_ GND GND VDD VDD _048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_47 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_133 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_3_166 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_3_177 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xhold6 net7 GND GND VDD VDD net27 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_3_Right_3 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_0_169 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_125 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_69 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk GND GND VDD VDD clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_2_209 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_15 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_088_ count\[1\] count\[2\] count\[3\] count\[0\] GND GND VDD VDD _047_ sky130_fd_sc_hd__or4b_1
XFILLER_3_189 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_48 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 _014_ GND GND VDD VDD net28 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_8_248 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_137 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_273 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_2_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_1_210 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_173 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_3_81 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_8_15 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_087_ _045_ _046_ _030_ GND GND VDD VDD _008_ sky130_fd_sc_hd__a21oi_1
Xhold8 net4 GND GND VDD VDD net29 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_113 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_49 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_91 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_1_233 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_1_222 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_9_141 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_130 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_9_185 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_15 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_086_ net1 _026_ _043_ GND GND VDD VDD _046_ sky130_fd_sc_hd__mux2_1
XFILLER_8_27 GND GND VDD VDD sky130_fd_sc_hd__fill_1
Xhold9 net9 GND GND VDD VDD net30 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_125 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_069_ net19 _032_ GND GND VDD VDD _034_ sky130_fd_sc_hd__or2_1
XFILLER_9_81 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_253 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_197 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_9_153 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_085_ count\[0\] count\[2\] count\[3\] count\[1\] GND GND VDD VDD _045_ sky130_fd_sc_hd__or4b_1
XFILLER_3_159 GND GND VDD VDD sky130_fd_sc_hd__fill_2
X_068_ net2 _029_ _032_ _033_ GND GND VDD VDD _002_ sky130_fd_sc_hd__and4_1
XFILLER_8_218 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_50 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_6_83 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_1_279 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_9_165 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_51 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_6_102 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_084_ _043_ _044_ _030_ GND GND VDD VDD _007_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_29 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_067_ net20 net21 count\[2\] GND GND VDD VDD _033_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_5_19 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_51 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_263 GND GND VDD VDD sky130_fd_sc_hd__fill_1
X_119_ clknet_1_1__leaf_clk net23 GND GND VDD VDD net8 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_285 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_1_225 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_7_3 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_9_111 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_6_114 GND GND VDD VDD sky130_fd_sc_hd__decap_8
X_083_ net1 _025_ _041_ GND GND VDD VDD _044_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_9_Left_19 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_3_139 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_97 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_53 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_066_ net20 net21 count\[2\] GND GND VDD VDD _032_ sky130_fd_sc_hd__nand3_2
XFILLER_2_183 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_0_109 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_52 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_253 GND GND VDD VDD sky130_fd_sc_hd__fill_2
X_118_ clknet_1_1__leaf_clk net28 GND GND VDD VDD net7 sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 net13 GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_6_41 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XFILLER_6_85 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_7 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_1_259 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_0_281 GND GND VDD VDD sky130_fd_sc_hd__decap_3
Xoutput3 net3 GND GND VDD VDD ADC0 sky130_fd_sc_hd__buf_2
X_082_ count\[2\] net19 net20 net21 GND GND VDD VDD _043_ sky130_fd_sc_hd__or4bb_1
X_065_ net20 net21 _031_ GND GND VDD VDD _001_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_195 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_9_85 GND GND VDD VDD sky130_fd_sc_hd__fill_2
XFILLER_9_52 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_9_41 GND GND VDD VDD sky130_fd_sc_hd__decap_6
X_117_ clknet_1_1__leaf_clk net34 GND GND VDD VDD net6 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_53 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_2 net13 GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_6_53 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xoutput4 net4 GND GND VDD VDD ADC1 sky130_fd_sc_hd__buf_2
XFILLER_9_113 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_10 GND GND VDD VDD sky130_fd_sc_hd__decap_3
X_081_ _041_ _042_ _030_ GND GND VDD VDD _006_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_149 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_3_108 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_2_130 GND GND VDD VDD sky130_fd_sc_hd__fill_1
X_064_ net20 net21 net2 GND GND VDD VDD _031_ sky130_fd_sc_hd__o21ai_1
X_116_ clknet_1_1__leaf_clk _012_ GND GND VDD VDD net5 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_54 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_233 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_4_214 VDD GND VDD GND sky130_ef_sc_hd__decap_12
XANTENNA_3 net13 GND GND VDD VDD sky130_fd_sc_hd__diode_2
XFILLER_6_65 VDD GND VDD GND sky130_ef_sc_hd__decap_12
Xoutput5 net5 GND GND VDD VDD ADC2 sky130_fd_sc_hd__buf_2
XFILLER_9_125 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_9_103 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_3_55 GND GND VDD VDD sky130_fd_sc_hd__fill_1
X_080_ net1 _024_ _039_ GND GND VDD VDD _042_ sky130_fd_sc_hd__mux2_1
XFILLER_6_139 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_65 GND VDD sky130_fd_sc_hd__tapvpwrvgnd_1
X_063_ net21 _030_ GND GND VDD VDD _000_ sky130_fd_sc_hd__nor2_1
XFILLER_2_197 VDD GND VDD GND sky130_ef_sc_hd__decap_12
X_115_ clknet_1_1__leaf_clk _011_ GND GND VDD VDD net4 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_223 GND GND VDD VDD sky130_fd_sc_hd__fill_1
XFILLER_7_245 GND GND VDD VDD sky130_fd_sc_hd__decap_8
XFILLER_4_226 GND GND VDD VDD sky130_fd_sc_hd__decap_6
XFILLER_4_248 GND GND VDD VDD sky130_fd_sc_hd__decap_4
XFILLER_3_281 GND GND VDD VDD sky130_fd_sc_hd__decap_3
XFILLER_6_77 GND GND VDD VDD sky130_fd_sc_hd__decap_6
Xoutput6 net6 GND GND VDD VDD ADC3 sky130_fd_sc_hd__buf_2
XFILLER_0_251 GND GND VDD VDD sky130_fd_sc_hd__fill_1
.ends

