magic
tech sky130A
timestamp 1759518789
<< nwell >>
rect -120 130 85 520
<< nmos >>
rect -50 -5 -35 95
<< pmos >>
rect -50 150 -35 250
<< ndiff >>
rect -100 80 -50 95
rect -100 10 -85 80
rect -65 10 -50 80
rect -100 -5 -50 10
rect -35 80 15 95
rect -35 10 -20 80
rect 0 10 15 80
rect -35 -5 15 10
<< pdiff >>
rect -100 235 -50 250
rect -100 165 -85 235
rect -65 165 -50 235
rect -100 150 -50 165
rect -35 235 15 250
rect -35 165 -20 235
rect 0 165 15 235
rect -35 150 15 165
<< ndiffc >>
rect -85 10 -65 80
rect -20 10 0 80
<< pdiffc >>
rect -85 165 -65 235
rect -20 165 0 235
<< psubdiff >>
rect 15 80 85 95
rect 15 10 30 80
rect 50 10 85 80
rect 15 -5 85 10
<< nsubdiff >>
rect 15 235 65 250
rect 15 165 30 235
rect 50 165 65 235
rect 15 150 65 165
<< psubdiffcont >>
rect 30 10 50 80
<< nsubdiffcont >>
rect 30 165 50 235
<< poly >>
rect -75 370 -35 380
rect -75 350 -65 370
rect -45 350 -35 370
rect -75 340 -35 350
rect -50 250 -35 340
rect -50 95 -35 150
rect -50 -20 -35 -5
<< polycont >>
rect -65 350 -45 370
<< locali >>
rect -120 435 85 455
rect -55 380 -35 435
rect -75 370 -35 380
rect -75 350 -65 370
rect -45 350 -35 370
rect -75 340 -35 350
rect -95 240 -75 245
rect -95 235 -55 240
rect -95 165 -85 235
rect -65 165 -55 235
rect -95 155 -55 165
rect -30 235 60 240
rect -30 165 -20 235
rect 0 165 30 235
rect 50 165 60 235
rect -30 155 60 165
rect -75 135 -55 155
rect 80 135 100 245
rect -75 115 100 135
rect -75 90 -55 115
rect -95 80 -55 90
rect -95 10 -85 80
rect -65 10 -55 80
rect -95 0 -55 10
rect -30 80 60 90
rect -30 10 -20 80
rect 0 10 30 80
rect 50 10 60 80
rect -30 0 60 10
<< viali >>
rect 30 165 50 235
rect 30 10 50 80
<< metal1 >>
rect -120 235 85 460
rect -120 165 30 235
rect 50 165 85 235
rect -120 150 85 165
rect -120 80 85 95
rect -120 10 30 80
rect 50 10 85 80
rect -120 -200 85 10
<< labels >>
rlabel locali -120 445 -120 445 7 A
port 0 w
rlabel locali 85 235 85 235 3 Y
port 1 e
rlabel metal1 -120 320 -120 320 7 VP
port 2 w
rlabel metal1 -120 -50 -120 -50 7 VN
port 3 w
<< end >>
