magic
tech sky130A
timestamp 1761856542
<< error_p >>
rect -390 -30 -365 270
rect -65 -30 -15 270
rect 285 -30 310 270
rect 610 -30 635 270
rect 935 -30 985 270
rect -470 -385 -420 -85
rect -120 -385 -70 -85
rect 230 -385 280 -85
rect 310 -385 360 -85
rect 660 -385 710 -85
rect 1010 -385 1060 -85
<< nmos >>
rect -365 -30 -65 270
rect -15 -30 285 270
rect 310 -30 610 270
rect 635 -30 935 270
rect -420 -385 -120 -85
rect -70 -385 230 -85
rect 360 -385 660 -85
rect 710 -385 1010 -85
<< ndiff >>
rect -390 -30 -365 270
rect -65 255 -15 270
rect -65 -15 -50 255
rect -30 -15 -15 255
rect -65 -30 -15 -15
rect 285 -30 310 270
rect 610 -30 635 270
rect 935 255 985 270
rect 935 -15 950 255
rect 970 -15 985 255
rect 935 -30 985 -15
rect -470 -100 -420 -85
rect -470 -370 -455 -100
rect -435 -370 -420 -100
rect -470 -385 -420 -370
rect -120 -100 -70 -85
rect -120 -370 -105 -100
rect -85 -370 -70 -100
rect -120 -385 -70 -370
rect 230 -100 280 -85
rect 230 -370 245 -100
rect 265 -370 280 -100
rect 230 -385 280 -370
rect 310 -100 360 -85
rect 310 -370 325 -100
rect 345 -370 360 -100
rect 310 -385 360 -370
rect 660 -100 710 -85
rect 660 -370 675 -100
rect 695 -370 710 -100
rect 660 -385 710 -370
rect 1010 -100 1060 -85
rect 1010 -370 1025 -100
rect 1045 -370 1060 -100
rect 1010 -385 1060 -370
<< ndiffc >>
rect -50 -15 -30 255
rect 950 -15 970 255
rect -455 -370 -435 -100
rect -105 -370 -85 -100
rect 245 -370 265 -100
rect 325 -370 345 -100
rect 675 -370 695 -100
rect 1025 -370 1045 -100
<< poly >>
rect -365 270 -65 285
rect -15 270 285 285
rect 310 270 610 285
rect 635 270 935 285
rect -365 -45 -65 -30
rect -15 -45 285 -30
rect 310 -45 610 -30
rect 635 -45 935 -30
rect -365 -70 -120 -45
rect -15 -70 230 -45
rect -420 -85 -120 -70
rect -70 -85 230 -70
rect 360 -70 610 -45
rect 710 -70 935 -45
rect 360 -85 660 -70
rect 710 -85 1010 -70
rect -420 -400 -120 -385
rect -70 -400 230 -385
rect 360 -400 660 -385
rect 710 -400 1010 -385
<< locali >>
rect -60 255 -20 265
rect -60 -15 -50 255
rect -30 -15 -20 255
rect -60 -25 -20 -15
rect 940 255 980 265
rect 940 -15 950 255
rect 970 -15 980 255
rect 940 -25 980 -15
rect -465 -100 -425 -90
rect -465 -370 -455 -100
rect -435 -370 -425 -100
rect -465 -400 -425 -370
rect -115 -100 -75 -90
rect -115 -370 -105 -100
rect -85 -370 -75 -100
rect -115 -380 -75 -370
rect 235 -100 275 -90
rect 235 -370 245 -100
rect 265 -370 275 -100
rect 235 -400 275 -370
rect -465 -420 275 -400
rect 315 -100 355 -90
rect 315 -370 325 -100
rect 345 -370 355 -100
rect 315 -400 355 -370
rect 665 -100 705 -90
rect 665 -370 675 -100
rect 695 -370 705 -100
rect 665 -380 705 -370
rect 1015 -100 1055 -90
rect 1015 -370 1025 -100
rect 1045 -370 1055 -100
rect 1015 -400 1055 -370
rect 315 -420 1055 -400
<< end >>
