magic
tech sky130A
timestamp 1762116719
<< nmos >>
rect 2600 7200 2800 8100
rect -200 6850 200 7150
rect 400 6850 800 7150
rect 900 7050 1100 7100
rect 1650 6250 1850 7150
rect 2100 6250 2300 7150
rect 2600 6250 2800 7150
rect -200 5900 200 6200
rect 400 5900 800 6200
rect 900 6100 1100 6150
rect 1650 5300 1850 6200
rect 2100 5300 2300 6200
rect 2600 5300 2800 6200
rect -200 4950 200 5250
rect 400 4950 800 5250
rect 900 5150 1100 5200
rect 1650 4350 1850 5250
rect 2100 4350 2300 5250
rect 2600 4350 2800 5250
rect -200 4000 200 4300
rect 400 4000 800 4300
rect 900 4200 1100 4250
rect 1650 3400 1850 4300
rect 2100 3400 2300 4300
rect 2600 3400 2800 4300
rect -200 3050 200 3350
rect 400 3050 800 3350
rect 900 3250 1100 3300
rect 1650 2450 1850 3350
rect 2100 2450 2300 3350
rect 2600 2450 2800 3350
rect -200 2100 200 2400
rect 400 2100 800 2400
rect 900 2300 1100 2350
rect 1650 1500 1850 2400
rect 2100 1500 2300 2400
rect 2600 1500 2800 2400
rect -200 1150 200 1450
rect 400 1150 800 1450
rect 900 1350 1100 1400
rect 2600 550 2800 1450
rect 2600 -400 2800 500
<< ndiff >>
rect 2350 8000 2600 8100
rect 2350 7300 2450 8000
rect 2500 7300 2600 8000
rect 2350 7200 2600 7300
rect 2800 8000 3050 8100
rect 2800 7300 2900 8000
rect 2950 7300 3050 8000
rect 2800 7200 3050 7300
rect -400 7050 -200 7150
rect -400 6950 -350 7050
rect -250 6950 -200 7050
rect -400 6850 -200 6950
rect 200 6850 400 7150
rect 800 7100 850 7150
rect 1400 7100 1650 7150
rect 800 7050 900 7100
rect 1100 7050 1650 7100
rect 800 6850 850 7050
rect 1400 6800 1500 7050
rect 1450 6750 1500 6800
rect 1400 6350 1500 6750
rect 1550 6350 1650 7050
rect 1400 6250 1650 6350
rect 1850 6600 2100 7150
rect 1850 6300 1950 6600
rect 2000 6300 2100 6600
rect 1850 6250 2100 6300
rect 2300 7050 2600 7150
rect 2300 6350 2450 7050
rect 2500 6350 2600 7050
rect 2300 6250 2600 6350
rect 2800 7050 3050 7150
rect 2800 6350 2900 7050
rect 2950 6350 3050 7050
rect 2800 6250 3050 6350
rect -400 6100 -200 6200
rect -400 6000 -350 6100
rect -250 6000 -200 6100
rect -400 5900 -200 6000
rect 200 5900 400 6200
rect 800 6150 850 6200
rect 1400 6150 1650 6200
rect 800 6100 900 6150
rect 1100 6100 1650 6150
rect 800 5900 850 6100
rect 1400 5850 1500 6100
rect 1450 5800 1500 5850
rect 1400 5400 1500 5800
rect 1550 5400 1650 6100
rect 1400 5300 1650 5400
rect 1850 5650 2100 6200
rect 1850 5350 1950 5650
rect 2000 5350 2100 5650
rect 1850 5300 2100 5350
rect 2300 6100 2600 6200
rect 2300 5400 2450 6100
rect 2500 5400 2600 6100
rect 2300 5300 2600 5400
rect 2800 6100 3050 6200
rect 2800 5400 2900 6100
rect 2950 5400 3050 6100
rect 2800 5300 3050 5400
rect -400 5150 -200 5250
rect -400 5050 -350 5150
rect -250 5050 -200 5150
rect -400 4950 -200 5050
rect 200 4950 400 5250
rect 800 5200 850 5250
rect 1400 5200 1650 5250
rect 800 5150 900 5200
rect 1100 5150 1650 5200
rect 800 4950 850 5150
rect 1400 4900 1500 5150
rect 1450 4850 1500 4900
rect 1400 4450 1500 4850
rect 1550 4450 1650 5150
rect 1400 4350 1650 4450
rect 1850 4700 2100 5250
rect 1850 4400 1950 4700
rect 2000 4400 2100 4700
rect 1850 4350 2100 4400
rect 2300 5150 2600 5250
rect 2300 4450 2450 5150
rect 2500 4450 2600 5150
rect 2300 4350 2600 4450
rect 2800 5150 3050 5250
rect 2800 4450 2900 5150
rect 2950 4450 3050 5150
rect 2800 4350 3050 4450
rect -400 4200 -200 4300
rect -400 4100 -350 4200
rect -250 4100 -200 4200
rect -400 4000 -200 4100
rect 200 4000 400 4300
rect 800 4250 850 4300
rect 1400 4250 1650 4300
rect 800 4200 900 4250
rect 1100 4200 1650 4250
rect 800 4000 850 4200
rect 1400 3950 1500 4200
rect 1450 3900 1500 3950
rect 1400 3500 1500 3900
rect 1550 3500 1650 4200
rect 1400 3400 1650 3500
rect 1850 3750 2100 4300
rect 1850 3450 1950 3750
rect 2000 3450 2100 3750
rect 1850 3400 2100 3450
rect 2300 4200 2600 4300
rect 2300 3500 2450 4200
rect 2500 3500 2600 4200
rect 2300 3400 2600 3500
rect 2800 4200 3050 4300
rect 2800 3500 2900 4200
rect 2950 3500 3050 4200
rect 2800 3400 3050 3500
rect -400 3250 -200 3350
rect -400 3150 -350 3250
rect -250 3150 -200 3250
rect -400 3050 -200 3150
rect 200 3050 400 3350
rect 800 3300 850 3350
rect 1400 3300 1650 3350
rect 800 3250 900 3300
rect 1100 3250 1650 3300
rect 800 3050 850 3250
rect 1400 3000 1500 3250
rect 1450 2950 1500 3000
rect 1400 2550 1500 2950
rect 1550 2550 1650 3250
rect 1400 2450 1650 2550
rect 1850 2800 2100 3350
rect 1850 2500 1950 2800
rect 2000 2500 2100 2800
rect 1850 2450 2100 2500
rect 2300 3250 2600 3350
rect 2300 2550 2450 3250
rect 2500 2550 2600 3250
rect 2300 2450 2600 2550
rect 2800 3250 3050 3350
rect 2800 2550 2900 3250
rect 2950 2550 3050 3250
rect 2800 2450 3050 2550
rect -400 2300 -200 2400
rect -400 2200 -350 2300
rect -250 2200 -200 2300
rect -400 2100 -200 2200
rect 200 2100 400 2400
rect 800 2350 850 2400
rect 1400 2350 1650 2400
rect 800 2300 900 2350
rect 1100 2300 1650 2350
rect 800 2100 850 2300
rect 1400 2050 1500 2300
rect 1450 2000 1500 2050
rect 1400 1600 1500 2000
rect 1550 1600 1650 2300
rect 1400 1500 1650 1600
rect 1850 1850 2100 2400
rect 1850 1550 1950 1850
rect 2000 1550 2100 1850
rect 1850 1500 2100 1550
rect 2300 2300 2600 2400
rect 2300 1600 2450 2300
rect 2500 1600 2600 2300
rect 2300 1500 2600 1600
rect 2800 2300 3050 2400
rect 2800 1600 2900 2300
rect 2950 1600 3050 2300
rect 2800 1500 3050 1600
rect -400 1350 -200 1450
rect -400 1250 -350 1350
rect -250 1250 -200 1350
rect -400 1150 -200 1250
rect 200 1150 400 1450
rect 800 1400 850 1450
rect 1400 1400 1600 1450
rect 800 1350 900 1400
rect 1100 1350 1600 1400
rect 800 1150 850 1350
rect 1400 1100 1500 1350
rect 1450 1050 1500 1100
rect 1400 650 1500 1050
rect 1550 650 1600 1350
rect 2350 1350 2600 1450
rect 1400 550 1600 650
rect 2350 650 2450 1350
rect 2500 650 2600 1350
rect 2350 550 2600 650
rect 2800 1350 3050 1450
rect 2800 650 2900 1350
rect 2950 650 3050 1350
rect 2800 550 3050 650
rect 2350 400 2600 500
rect 2350 -300 2450 400
rect 2500 -300 2600 400
rect 2350 -400 2600 -300
rect 2800 400 3050 500
rect 2800 -300 2900 400
rect 2950 -300 3050 400
rect 2800 -400 3050 -300
<< ndiffc >>
rect 2450 7300 2500 8000
rect 2900 7300 2950 8000
rect -350 6950 -250 7050
rect 1500 6350 1550 7050
rect 1950 6300 2000 6600
rect 2450 6350 2500 7050
rect 2900 6350 2950 7050
rect -350 6000 -250 6100
rect 1500 5400 1550 6100
rect 1950 5350 2000 5650
rect 2450 5400 2500 6100
rect 2900 5400 2950 6100
rect -350 5050 -250 5150
rect 1500 4450 1550 5150
rect 1950 4400 2000 4700
rect 2450 4450 2500 5150
rect 2900 4450 2950 5150
rect -350 4100 -250 4200
rect 1500 3500 1550 4200
rect 1950 3450 2000 3750
rect 2450 3500 2500 4200
rect 2900 3500 2950 4200
rect -350 3150 -250 3250
rect 1500 2550 1550 3250
rect 1950 2500 2000 2800
rect 2450 2550 2500 3250
rect 2900 2550 2950 3250
rect -350 2200 -250 2300
rect 1500 1600 1550 2300
rect 1950 1550 2000 1850
rect 2450 1600 2500 2300
rect 2900 1600 2950 2300
rect -350 1250 -250 1350
rect 1500 650 1550 1350
rect 2450 650 2500 1350
rect 2900 650 2950 1350
rect 2450 -300 2500 400
rect 2900 -300 2950 400
<< psubdiff >>
rect 3050 8000 3300 8100
rect 3050 7300 3150 8000
rect 3200 7300 3300 8000
rect 3050 7200 3300 7300
rect -600 7050 -400 7150
rect -600 6950 -550 7050
rect -450 6950 -400 7050
rect -600 6850 -400 6950
rect 1150 6650 1400 6750
rect 1150 6350 1250 6650
rect 1300 6350 1400 6650
rect 1150 6250 1400 6350
rect -600 6100 -400 6200
rect -600 6000 -550 6100
rect -450 6000 -400 6100
rect -600 5900 -400 6000
rect 1150 5700 1400 5800
rect 1150 5400 1250 5700
rect 1300 5400 1400 5700
rect 1150 5300 1400 5400
rect 3050 6100 3300 6200
rect 3050 5400 3150 6100
rect 3200 5400 3300 6100
rect 3050 5300 3300 5400
rect -600 5150 -400 5250
rect -600 5050 -550 5150
rect -450 5050 -400 5150
rect -600 4950 -400 5050
rect 1150 4750 1400 4850
rect 1150 4450 1250 4750
rect 1300 4450 1400 4750
rect 1150 4350 1400 4450
rect -600 4200 -400 4300
rect -600 4100 -550 4200
rect -450 4100 -400 4200
rect -600 4000 -400 4100
rect 1150 3800 1400 3900
rect 1150 3500 1250 3800
rect 1300 3500 1400 3800
rect 1150 3400 1400 3500
rect 3050 4200 3300 4300
rect 3050 3500 3150 4200
rect 3200 3500 3300 4200
rect 3050 3400 3300 3500
rect -600 3250 -400 3350
rect -600 3150 -550 3250
rect -450 3150 -400 3250
rect -600 3050 -400 3150
rect 1150 2850 1400 2950
rect 1150 2550 1250 2850
rect 1300 2550 1400 2850
rect 1150 2450 1400 2550
rect -600 2300 -400 2400
rect -600 2200 -550 2300
rect -450 2200 -400 2300
rect -600 2100 -400 2200
rect 1150 1900 1400 2000
rect 1150 1600 1250 1900
rect 1300 1600 1400 1900
rect 1150 1500 1400 1600
rect 3050 2300 3300 2400
rect 3050 1600 3150 2300
rect 3200 1600 3300 2300
rect 3050 1500 3300 1600
rect -600 1350 -400 1450
rect -600 1250 -550 1350
rect -450 1250 -400 1350
rect -600 1150 -400 1250
rect 1150 950 1400 1050
rect 1150 650 1250 950
rect 1300 650 1400 950
rect 1150 550 1400 650
rect 3050 400 3300 500
rect 3050 -300 3150 400
rect 3200 -300 3300 400
rect 3050 -400 3300 -300
<< psubdiffcont >>
rect 3150 7300 3200 8000
rect -550 6950 -450 7050
rect 1250 6350 1300 6650
rect -550 6000 -450 6100
rect 1250 5400 1300 5700
rect 3150 5400 3200 6100
rect -550 5050 -450 5150
rect 1250 4450 1300 4750
rect -550 4100 -450 4200
rect 1250 3500 1300 3800
rect 3150 3500 3200 4200
rect -550 3150 -450 3250
rect 1250 2550 1300 2850
rect -550 2200 -450 2300
rect 1250 1600 1300 1900
rect 3150 1600 3200 2300
rect -550 1250 -450 1350
rect 1250 650 1300 950
rect 3150 -300 3200 400
<< poly >>
rect 1650 8300 1850 8350
rect -200 8250 200 8300
rect -200 8150 -150 8250
rect 150 8150 200 8250
rect -200 7150 200 8150
rect 400 8250 800 8300
rect 400 8150 450 8250
rect 750 8150 800 8250
rect 400 7150 800 8150
rect 1650 8200 1700 8300
rect 1800 8200 1850 8300
rect 1650 7150 1850 8200
rect 2100 8300 2300 8350
rect 2100 8200 2150 8300
rect 2250 8200 2300 8300
rect 2100 7150 2300 8200
rect 2600 8300 2800 8350
rect 2600 8200 2650 8300
rect 2750 8200 2800 8300
rect 2600 8100 2800 8200
rect 2600 7150 2800 7200
rect 900 7100 1100 7150
rect -200 6200 200 6850
rect 400 6200 800 6850
rect 900 6400 1100 7050
rect 900 6300 950 6400
rect 1050 6300 1100 6400
rect 900 6250 1100 6300
rect 1650 6200 1850 6250
rect 2100 6200 2300 6250
rect 2600 6200 2800 6250
rect 900 6150 1100 6200
rect -200 5250 200 5900
rect 400 5250 800 5900
rect 900 5450 1100 6100
rect 900 5350 950 5450
rect 1050 5350 1100 5450
rect 900 5300 1100 5350
rect 1650 5250 1850 5300
rect 2100 5250 2300 5300
rect 2600 5250 2800 5300
rect 900 5200 1100 5250
rect -200 4300 200 4950
rect 400 4300 800 4950
rect 900 4500 1100 5150
rect 900 4400 950 4500
rect 1050 4400 1100 4500
rect 900 4350 1100 4400
rect 1650 4300 1850 4350
rect 2100 4300 2300 4350
rect 2600 4300 2800 4350
rect 900 4250 1100 4300
rect -200 3350 200 4000
rect 400 3350 800 4000
rect 900 3550 1100 4200
rect 900 3450 950 3550
rect 1050 3450 1100 3550
rect 900 3400 1100 3450
rect 1650 3350 1850 3400
rect 2100 3350 2300 3400
rect 2600 3350 2800 3400
rect 900 3300 1100 3350
rect -200 2400 200 3050
rect 400 2400 800 3050
rect 900 2600 1100 3250
rect 900 2500 950 2600
rect 1050 2500 1100 2600
rect 900 2450 1100 2500
rect 1650 2400 1850 2450
rect 2100 2400 2300 2450
rect 2600 2400 2800 2450
rect 900 2350 1100 2400
rect -200 1450 200 2100
rect 400 1450 800 2100
rect 900 1650 1100 2300
rect 900 1550 950 1650
rect 1050 1550 1100 1650
rect 900 1500 1100 1550
rect 900 1400 1100 1450
rect -200 1100 200 1150
rect 400 1100 800 1150
rect 900 700 1100 1350
rect 900 600 950 700
rect 1050 600 1100 700
rect 900 550 1100 600
rect 1650 950 1850 1500
rect 2100 950 2300 1500
rect 2600 1450 2800 1500
rect 2600 500 2800 550
rect 2600 -550 2800 -400
<< polycont >>
rect -150 8150 150 8250
rect 450 8150 750 8250
rect 1700 8200 1800 8300
rect 2150 8200 2250 8300
rect 2650 8200 2750 8300
rect 950 6300 1050 6400
rect 950 5350 1050 5450
rect 950 4400 1050 4500
rect 950 3450 1050 3550
rect 950 2500 1050 2600
rect 950 1550 1050 1650
rect 950 600 1050 700
<< locali >>
rect -650 8700 1650 8850
rect -650 8500 800 8650
rect -650 8300 200 8450
rect -200 8250 200 8300
rect -200 8150 -150 8250
rect 150 8150 200 8250
rect -200 8100 200 8150
rect 400 8250 800 8500
rect 400 8150 450 8250
rect 750 8150 800 8250
rect 1450 8350 1650 8700
rect 1450 8300 2800 8350
rect 1450 8200 1700 8300
rect 1800 8200 2150 8300
rect 2250 8200 2650 8300
rect 2750 8200 2800 8300
rect 1450 8150 2800 8200
rect 400 8100 800 8150
rect 2400 8000 2550 8050
rect 2400 7300 2450 8000
rect 2500 7300 2550 8000
rect 2400 7100 2550 7300
rect -550 7050 -250 7100
rect -450 6950 -350 7050
rect -550 6900 -250 6950
rect -400 6850 -250 6900
rect 1450 7050 2550 7100
rect 1450 6700 1500 7050
rect 1200 6650 1350 6700
rect -650 6400 1100 6450
rect -650 6300 950 6400
rect 1050 6300 1100 6400
rect 1200 6350 1250 6650
rect 1300 6350 1350 6650
rect 1200 6300 1350 6350
rect 1400 6350 1500 6700
rect 1550 6700 2450 7050
rect 1550 6350 1600 6700
rect 1400 6300 1600 6350
rect 1900 6600 2050 6650
rect 1900 6300 1950 6600
rect 2000 6300 2050 6600
rect 2400 6350 2450 6700
rect 2500 6350 2550 7050
rect 2400 6300 2550 6350
rect 2850 8000 3050 8050
rect 2850 7300 2900 8000
rect 2950 7300 3050 8000
rect 2850 7250 3050 7300
rect 3100 8000 3250 8050
rect 3100 7300 3150 8000
rect 3200 7300 3250 8000
rect 3100 7250 3250 7300
rect 2850 7050 3000 7250
rect 2850 6350 2900 7050
rect 2950 6350 3000 7050
rect -650 6250 1100 6300
rect -400 6150 -250 6200
rect 1900 6150 2050 6300
rect 2850 6150 3000 6350
rect -550 6100 -250 6150
rect -450 6000 -350 6100
rect -550 5950 -250 6000
rect -400 5900 -250 5950
rect 1450 6100 2550 6150
rect 1200 5700 1350 5750
rect -650 5450 1100 5500
rect -650 5350 950 5450
rect 1050 5350 1100 5450
rect 1200 5400 1250 5700
rect 1300 5400 1350 5700
rect 1200 5350 1350 5400
rect 1450 5400 1500 6100
rect 1550 5750 2450 6100
rect 1550 5400 1600 5750
rect 1450 5350 1600 5400
rect 1900 5650 2050 5700
rect 1900 5350 1950 5650
rect 2000 5350 2050 5650
rect 2400 5400 2450 5750
rect 2500 5400 2550 6100
rect 2400 5350 2550 5400
rect 2850 6100 3050 6150
rect 2850 5400 2900 6100
rect 2950 5400 3050 6100
rect 2850 5350 3050 5400
rect 3100 6100 3250 6150
rect 3100 5400 3150 6100
rect 3200 5400 3250 6100
rect 3100 5350 3250 5400
rect -650 5300 1100 5350
rect -400 5200 -250 5250
rect 1900 5200 2050 5350
rect -550 5150 -250 5200
rect -450 5050 -350 5150
rect -550 5000 -250 5050
rect -400 4950 -250 5000
rect 1450 5150 2550 5200
rect 1200 4750 1350 4800
rect -650 4500 1100 4550
rect -650 4400 950 4500
rect 1050 4400 1100 4500
rect 1200 4450 1250 4750
rect 1300 4450 1350 4750
rect 1200 4400 1350 4450
rect 1450 4450 1500 5150
rect 1550 4800 2450 5150
rect 1550 4450 1600 4800
rect 1450 4400 1600 4450
rect 1900 4700 2050 4750
rect 1900 4400 1950 4700
rect 2000 4400 2050 4700
rect 2400 4450 2450 4800
rect 2500 4450 2550 5150
rect 2400 4400 2550 4450
rect 2850 5150 3000 5350
rect 2850 4450 2900 5150
rect 2950 4450 3000 5150
rect -650 4350 1100 4400
rect -400 4250 -250 4300
rect 1900 4250 2050 4400
rect 2850 4250 3000 4450
rect -550 4200 -250 4250
rect -450 4100 -350 4200
rect -550 4050 -250 4100
rect -400 4000 -250 4050
rect 1450 4200 2550 4250
rect 1200 3800 1350 3850
rect -650 3550 1100 3600
rect -650 3450 950 3550
rect 1050 3450 1100 3550
rect 1200 3500 1250 3800
rect 1300 3500 1350 3800
rect 1200 3450 1350 3500
rect 1450 3500 1500 4200
rect 1550 3850 2450 4200
rect 1550 3500 1600 3850
rect 1450 3450 1600 3500
rect 1900 3750 2050 3800
rect 1900 3450 1950 3750
rect 2000 3450 2050 3750
rect 2400 3500 2450 3850
rect 2500 3500 2550 4200
rect 2400 3450 2550 3500
rect 2850 4200 3050 4250
rect 2850 3500 2900 4200
rect 2950 3500 3050 4200
rect 2850 3450 3050 3500
rect 3100 4200 3250 4250
rect 3100 3500 3150 4200
rect 3200 3500 3250 4200
rect 3100 3450 3250 3500
rect -650 3400 1100 3450
rect -400 3300 -250 3350
rect 1900 3300 2050 3450
rect -550 3250 -250 3300
rect -450 3150 -350 3250
rect -550 3100 -250 3150
rect -400 3050 -250 3100
rect 1450 3250 2550 3300
rect 1200 2850 1350 2900
rect -650 2600 1100 2650
rect -650 2500 950 2600
rect 1050 2500 1100 2600
rect 1200 2550 1250 2850
rect 1300 2550 1350 2850
rect 1200 2500 1350 2550
rect 1450 2550 1500 3250
rect 1550 2900 2450 3250
rect 1550 2550 1600 2900
rect 1450 2500 1600 2550
rect 1900 2800 2050 2850
rect 1900 2500 1950 2800
rect 2000 2500 2050 2800
rect 2400 2550 2450 2900
rect 2500 2550 2550 3250
rect 2400 2500 2550 2550
rect 2850 3250 3000 3450
rect 2850 2550 2900 3250
rect 2950 2550 3000 3250
rect -650 2450 1100 2500
rect -400 2350 -250 2400
rect 1900 2350 2050 2500
rect 2850 2350 3000 2550
rect -550 2300 -250 2350
rect -450 2200 -350 2300
rect -550 2150 -250 2200
rect -400 2100 -250 2150
rect 1450 2300 2550 2350
rect 1200 1900 1350 1950
rect -650 1650 1100 1700
rect -650 1550 950 1650
rect 1050 1550 1100 1650
rect 1200 1600 1250 1900
rect 1300 1600 1350 1900
rect 1200 1550 1350 1600
rect 1450 1600 1500 2300
rect 1550 1950 2450 2300
rect 1550 1600 1600 1950
rect 1450 1550 1600 1600
rect 1900 1850 2050 1900
rect 1900 1550 1950 1850
rect 2000 1550 2050 1850
rect 2400 1600 2450 1950
rect 2500 1600 2550 2300
rect 2400 1550 2550 1600
rect 2850 2300 3050 2350
rect 2850 1600 2900 2300
rect 2950 1600 3050 2300
rect 2850 1550 3050 1600
rect 3100 2300 3250 2350
rect 3100 1600 3150 2300
rect 3200 1600 3250 2300
rect 3100 1550 3250 1600
rect -650 1500 1100 1550
rect -400 1400 -250 1450
rect 1900 1400 2050 1550
rect -550 1350 -250 1400
rect -450 1250 -350 1350
rect -550 1200 -250 1250
rect 1450 1350 2550 1400
rect 1200 950 1350 1000
rect -650 700 1100 750
rect -650 600 950 700
rect 1050 600 1100 700
rect 1200 650 1250 950
rect 1300 650 1350 950
rect 1200 600 1350 650
rect 1450 650 1500 1350
rect 1550 1000 2450 1350
rect 1550 650 1600 1000
rect 1450 600 1600 650
rect 2400 650 2450 1000
rect 2500 650 2550 1350
rect -650 550 1100 600
rect 2400 400 2550 650
rect 2400 -300 2450 400
rect 2500 -300 2550 400
rect 2400 -350 2550 -300
rect 2850 1350 3000 1400
rect 2850 650 2900 1350
rect 2950 650 3000 1350
rect 2850 400 3000 650
rect 2850 -300 2900 400
rect 2950 -300 3000 400
rect 2850 -450 3000 -300
rect 3100 400 3250 450
rect 3100 -300 3150 400
rect 3200 -300 3250 400
rect 3100 -350 3250 -300
rect 2850 -600 3350 -450
<< viali >>
rect -350 6950 -250 7050
rect 2900 7300 2950 8000
rect 2900 6350 2950 7050
rect -350 6000 -250 6100
rect 2900 5400 2950 6100
rect -350 5050 -250 5150
rect 2900 4450 2950 5150
rect -350 4100 -250 4200
rect 2900 3500 2950 4200
rect -350 3150 -250 3250
rect 2900 2550 2950 3250
rect -350 2200 -250 2300
rect 2900 1600 2950 2300
rect -350 1250 -250 1350
<< metal1 >>
rect -650 8000 3300 8100
rect -650 7300 2900 8000
rect 2950 7300 3300 8000
rect -650 7200 3300 7300
rect -550 7050 -200 7100
rect -550 6950 -350 7050
rect -250 6950 -200 7050
rect -550 6100 -200 6950
rect -550 6000 -350 6100
rect -250 6000 -200 6100
rect -550 5150 -200 6000
rect -550 5050 -350 5150
rect -250 5050 -200 5150
rect -550 4200 -200 5050
rect -550 4100 -350 4200
rect -250 4100 -200 4200
rect -550 3250 -200 4100
rect -550 3150 -350 3250
rect -250 3150 -200 3250
rect -550 2300 -200 3150
rect -550 2200 -350 2300
rect -250 2200 -200 2300
rect -550 1350 -200 2200
rect 2850 7050 3250 7200
rect 2850 6350 2900 7050
rect 2950 6350 3250 7050
rect 2850 6100 3250 6350
rect 2850 5400 2900 6100
rect 2950 5400 3250 6100
rect 2850 5150 3250 5400
rect 2850 4450 2900 5150
rect 2950 4450 3250 5150
rect 2850 4200 3250 4450
rect 2850 3500 2900 4200
rect 2950 3500 3250 4200
rect 2850 3250 3250 3500
rect 2850 2550 2900 3250
rect 2950 2550 3250 3250
rect 2850 2300 3250 2550
rect 2850 1600 2900 2300
rect 2950 1600 3250 2300
rect 2850 1500 3250 1600
rect -550 1250 -350 1350
rect -250 1250 -200 1350
rect -550 500 -200 1250
rect -650 -400 3350 500
<< labels >>
rlabel locali 3350 -550 3350 -550 3 Iout
port 1 e
rlabel locali -650 650 -650 650 3 D6
port 2 e
rlabel locali -650 1600 -650 1600 3 D5
port 3 e
rlabel locali -650 2550 -650 2550 3 D4
port 4 e
rlabel locali -650 3500 -650 3500 3 D3
port 5 e
rlabel locali -650 4450 -650 4450 3 D2
port 6 e
rlabel locali -650 5400 -650 5400 3 D1
port 7 e
rlabel locali -650 6350 -650 6350 3 D0
port 8 e
rlabel locali -650 8600 -650 8600 3 Vc
port 9 e
rlabel locali -650 8800 -650 8800 3 Vg
port 10 e
rlabel metal1 -650 50 -650 50 3 GND
port 11 e
rlabel locali -650 8400 -650 8400 3 Vbn
port 12 e
rlabel metal1 -650 7650 -650 7650 3 VDD
port 13 e
<< end >>
