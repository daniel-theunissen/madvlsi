magic
tech sky130A
timestamp 1759703914
<< nwell >>
rect -205 310 165 700
<< nmos >>
rect -105 175 -90 275
rect -65 175 -50 275
rect 0 175 45 275
rect 100 175 115 275
rect -105 -20 -90 80
rect -65 -20 -50 80
rect 0 -20 45 80
rect 100 -20 115 80
<< pmos >>
rect -125 540 -80 640
rect -30 540 -15 640
rect 35 540 50 640
rect 75 540 90 640
rect -125 330 -80 430
rect -30 330 -15 430
rect 35 330 50 430
rect 75 330 90 430
<< ndiff >>
rect -155 260 -105 275
rect -155 240 -140 260
rect -120 240 -105 260
rect -155 175 -105 240
rect -90 175 -65 275
rect -50 260 0 275
rect -50 190 -35 260
rect -15 190 0 260
rect -50 175 0 190
rect 45 260 100 275
rect 45 190 65 260
rect 85 190 100 260
rect 45 175 100 190
rect 115 260 165 275
rect 115 190 130 260
rect 150 190 165 260
rect 115 175 165 190
rect -155 15 -105 80
rect -155 -5 -140 15
rect -120 -5 -105 15
rect -155 -20 -105 -5
rect -90 -20 -65 80
rect -50 65 0 80
rect -50 -5 -35 65
rect -15 -5 0 65
rect -50 -20 0 -5
rect 45 65 100 80
rect 45 -5 65 65
rect 85 -5 100 65
rect 45 -20 100 -5
rect 115 65 165 80
rect 115 -5 130 65
rect 150 -5 165 65
rect 115 -20 165 -5
<< pdiff >>
rect -180 625 -125 640
rect -180 555 -165 625
rect -145 555 -125 625
rect -180 540 -125 555
rect -80 625 -30 640
rect -80 555 -65 625
rect -45 555 -30 625
rect -80 540 -30 555
rect -15 625 35 640
rect -15 555 0 625
rect 20 555 35 625
rect -15 540 35 555
rect 50 540 75 640
rect 90 625 140 640
rect 90 555 105 625
rect 125 555 140 625
rect 90 540 140 555
rect -175 415 -125 430
rect -175 345 -160 415
rect -140 345 -125 415
rect -175 330 -125 345
rect -80 415 -30 430
rect -80 345 -65 415
rect -45 345 -30 415
rect -80 330 -30 345
rect -15 415 35 430
rect -15 345 0 415
rect 20 345 35 415
rect -15 330 35 345
rect 50 330 75 430
rect 90 415 140 430
rect 90 345 105 415
rect 125 345 140 415
rect 90 330 140 345
<< ndiffc >>
rect -140 240 -120 260
rect -35 190 -15 260
rect 65 190 85 260
rect 130 190 150 260
rect -140 -5 -120 15
rect -35 -5 -15 65
rect 65 -5 85 65
rect 130 -5 150 65
<< pdiffc >>
rect -165 555 -145 625
rect -65 555 -45 625
rect 0 555 20 625
rect 105 555 125 625
rect -160 345 -140 415
rect -65 345 -45 415
rect 0 345 20 415
rect 105 345 125 415
<< psubdiff >>
rect -205 260 -155 275
rect -205 190 -190 260
rect -170 190 -155 260
rect -205 175 -155 190
rect -205 65 -155 80
rect -205 -5 -190 65
rect -170 -5 -155 65
rect -205 -20 -155 -5
<< nsubdiff >>
rect -185 495 -135 510
rect -185 475 -170 495
rect -150 475 -135 495
rect -185 460 -135 475
<< psubdiffcont >>
rect -190 190 -170 260
rect -190 -5 -170 65
<< nsubdiffcont >>
rect -170 475 -150 495
<< poly >>
rect -55 685 -15 695
rect -55 665 -45 685
rect -25 665 -15 685
rect -55 655 -15 665
rect 75 685 115 695
rect 75 665 85 685
rect 105 665 115 685
rect 75 655 115 665
rect -125 640 -80 655
rect -30 640 -15 655
rect 35 640 50 655
rect 75 640 90 655
rect -125 430 -80 540
rect -30 525 -15 540
rect -55 475 -15 485
rect -55 455 -45 475
rect -25 455 -15 475
rect -55 445 -15 455
rect -30 430 -15 445
rect 35 430 50 540
rect 75 525 90 540
rect 95 475 135 485
rect 95 455 105 475
rect 125 455 135 475
rect 75 445 135 455
rect 75 440 110 445
rect 75 430 90 440
rect -125 315 -80 330
rect -30 320 -15 330
rect -105 275 -90 315
rect -40 305 -15 320
rect 35 310 50 330
rect -40 300 -25 305
rect -65 285 -25 300
rect 30 290 50 310
rect 75 320 90 330
rect 75 305 115 320
rect -65 275 -50 285
rect 0 275 45 290
rect 100 275 115 305
rect -105 80 -90 175
rect -65 160 -50 175
rect -65 150 -25 160
rect -65 130 -55 150
rect -35 130 -25 150
rect -65 120 -25 130
rect -65 80 -50 95
rect 0 80 45 175
rect 100 160 115 175
rect 75 150 115 160
rect 75 130 85 150
rect 105 130 115 150
rect 75 120 115 130
rect 100 80 115 95
rect -105 -30 -90 -20
rect -130 -45 -90 -30
rect -130 -95 -115 -45
rect -65 -70 -50 -20
rect 0 -35 45 -20
rect 100 -35 115 -20
rect -155 -105 -115 -95
rect -155 -125 -145 -105
rect -125 -125 -115 -105
rect -90 -80 -50 -70
rect -90 -100 -80 -80
rect -60 -100 -50 -80
rect 30 -95 45 -35
rect 75 -45 115 -35
rect 75 -65 85 -45
rect 105 -65 115 -45
rect 75 -75 115 -65
rect -90 -110 -50 -100
rect 15 -105 55 -95
rect -155 -135 -115 -125
rect 15 -125 25 -105
rect 45 -125 55 -105
rect 15 -135 55 -125
<< polycont >>
rect -45 665 -25 685
rect 85 665 105 685
rect -45 455 -25 475
rect 105 455 125 475
rect -55 130 -35 150
rect 85 130 105 150
rect -145 -125 -125 -105
rect -80 -100 -60 -80
rect 85 -65 105 -45
rect 25 -125 45 -105
<< locali >>
rect -55 685 -15 695
rect -55 675 -45 685
rect -115 665 -45 675
rect -25 665 -15 685
rect 75 685 115 695
rect 75 675 85 685
rect -115 655 -15 665
rect 55 665 85 675
rect 105 665 115 685
rect 55 655 115 665
rect -205 625 -135 635
rect -205 615 -165 625
rect -175 555 -165 615
rect -145 555 -135 625
rect -175 545 -135 555
rect -180 495 -140 505
rect -180 475 -170 495
rect -150 475 -140 495
rect -180 465 -140 475
rect -115 455 -95 655
rect -75 625 -35 635
rect -75 555 -65 625
rect -45 555 -35 625
rect -75 545 -35 555
rect -10 625 30 635
rect -10 555 0 625
rect 20 555 30 625
rect -10 545 30 555
rect -55 485 -35 545
rect -55 475 -15 485
rect -55 455 -45 475
rect -25 455 -15 475
rect -115 445 -90 455
rect -55 445 -15 455
rect -110 425 -90 445
rect 10 425 30 545
rect -205 415 -130 425
rect -205 405 -160 415
rect -170 345 -160 405
rect -140 345 -130 415
rect -110 415 -35 425
rect -110 405 -65 415
rect -170 335 -130 345
rect -75 345 -65 405
rect -45 345 -35 415
rect -75 335 -35 345
rect -10 415 30 425
rect -10 345 0 415
rect 20 345 30 415
rect 55 425 75 655
rect 145 635 165 700
rect 95 625 165 635
rect 95 555 105 625
rect 125 615 165 625
rect 125 555 135 615
rect 95 545 135 555
rect 95 485 115 545
rect 95 475 135 485
rect 95 455 105 475
rect 125 455 135 475
rect 95 445 135 455
rect 55 415 165 425
rect 55 405 105 415
rect 95 355 105 405
rect -10 335 30 345
rect 85 345 105 355
rect 125 405 165 415
rect 125 345 135 405
rect 85 335 135 345
rect -55 320 -35 335
rect 85 330 105 335
rect -55 305 -25 320
rect -45 270 -25 305
rect 75 315 105 330
rect 75 270 95 315
rect -205 260 -110 270
rect -205 190 -190 260
rect -170 240 -140 260
rect -120 240 -110 260
rect -170 230 -110 240
rect -45 260 -5 270
rect -170 190 -130 230
rect -45 200 -35 260
rect -205 180 -130 190
rect -150 75 -130 180
rect -110 190 -35 200
rect -15 190 -5 260
rect 55 260 95 270
rect 55 200 65 260
rect -110 180 -5 190
rect 15 190 65 200
rect 85 190 95 260
rect 15 180 95 190
rect 120 260 165 270
rect 120 190 130 260
rect 150 190 165 260
rect 120 180 165 190
rect -110 100 -85 180
rect -65 150 -25 160
rect -65 130 -55 150
rect -35 130 -25 150
rect -65 120 -25 130
rect -110 80 -70 100
rect -205 65 -130 75
rect -205 -5 -190 65
rect -170 25 -130 65
rect -170 15 -110 25
rect -170 -5 -140 15
rect -120 -5 -110 15
rect -205 -15 -110 -5
rect -90 -70 -70 80
rect -45 75 -25 120
rect -45 65 -5 75
rect -45 -5 -35 65
rect -15 -5 -5 65
rect -45 -15 -5 -5
rect 15 -35 35 180
rect 75 150 115 160
rect 75 130 85 150
rect 105 130 115 150
rect 75 120 115 130
rect 75 75 95 120
rect 140 75 160 180
rect 55 65 95 75
rect 55 -5 65 65
rect 85 -5 95 65
rect 55 -15 95 -5
rect 120 65 165 75
rect 120 -5 130 65
rect 150 -5 165 65
rect 120 -15 165 -5
rect 15 -45 115 -35
rect 15 -55 85 -45
rect 75 -65 85 -55
rect 105 -65 115 -45
rect -90 -80 -50 -70
rect 75 -75 115 -65
rect -155 -105 -115 -95
rect -155 -125 -145 -105
rect -125 -125 -115 -105
rect -90 -100 -80 -80
rect -60 -100 -50 -80
rect -90 -110 -50 -100
rect 15 -105 55 -95
rect -155 -135 -115 -125
rect 15 -125 25 -105
rect 45 -125 55 -105
rect 15 -135 55 -125
<< viali >>
rect -170 475 -150 495
rect 0 555 20 625
rect 0 345 20 415
rect -190 190 -170 260
rect -140 240 -120 260
rect 130 190 150 260
rect -190 -5 -170 65
rect -140 -5 -120 15
rect 130 -5 150 65
rect -145 -125 -125 -105
rect 25 -125 45 -105
<< metal1 >>
rect -205 625 165 640
rect -205 555 0 625
rect 20 555 165 625
rect -205 495 165 555
rect -205 475 -170 495
rect -150 475 165 495
rect -205 415 165 475
rect -205 345 0 415
rect 20 345 165 415
rect -205 330 165 345
rect -205 260 165 275
rect -205 190 -190 260
rect -170 240 -140 260
rect -120 240 130 260
rect -170 190 130 240
rect 150 190 165 260
rect -205 65 165 190
rect -205 -5 -190 65
rect -170 15 130 65
rect -170 -5 -140 15
rect -120 -5 130 15
rect 150 -5 165 65
rect -205 -20 165 -5
rect -205 -105 165 -95
rect -205 -125 -145 -105
rect -125 -125 25 -105
rect 45 -125 165 -105
rect -205 -135 165 -125
<< labels >>
rlabel metal1 -205 -115 -205 -115 7 clk
port 0 w
rlabel locali 165 625 165 625 3 Q
port 3 e
rlabel locali 165 415 165 415 3 Qn
port 4 e
rlabel metal1 -205 485 -205 485 7 VP
port 5 w
rlabel metal1 -205 125 -205 125 7 VN
port 6 w
rlabel locali -205 625 -205 625 7 D
port 1 w
rlabel locali -205 415 -205 415 7 Dn
port 2 w
<< end >>
